magic
tech scmos
timestamp 1638815411
<< nwell >>
rect -268 191 622 218
rect -343 123 667 150
rect -290 4 651 31
<< ntransistor >>
rect -257 165 -255 169
rect -247 165 -245 169
rect -230 165 -228 169
rect -220 165 -218 169
rect -210 165 -208 169
rect -200 165 -198 169
rect -184 165 -182 169
rect -174 165 -172 169
rect -164 165 -162 169
rect -148 165 -146 169
rect -138 165 -136 169
rect -121 165 -119 169
rect -111 165 -109 169
rect -101 165 -99 169
rect -91 165 -89 169
rect -75 165 -73 169
rect -65 165 -63 169
rect -55 165 -53 169
rect -29 165 -27 169
rect -19 165 -17 169
rect -2 165 0 169
rect 8 165 10 169
rect 18 165 20 169
rect 28 165 30 169
rect 44 165 46 169
rect 54 165 56 169
rect 64 165 66 169
rect 80 165 82 169
rect 90 165 92 169
rect 107 165 109 169
rect 117 165 119 169
rect 127 165 129 169
rect 137 165 139 169
rect 153 165 155 169
rect 163 165 165 169
rect 173 165 175 169
rect 189 165 191 169
rect 199 165 201 169
rect 216 165 218 169
rect 226 165 228 169
rect 236 165 238 169
rect 246 165 248 169
rect 262 165 264 169
rect 272 165 274 169
rect 282 165 284 169
rect 298 165 300 169
rect 308 165 310 169
rect 325 165 327 169
rect 335 165 337 169
rect 345 165 347 169
rect 355 165 357 169
rect 371 165 373 169
rect 381 165 383 169
rect 391 165 393 169
rect 407 165 409 169
rect 417 165 419 169
rect 434 165 436 169
rect 444 165 446 169
rect 454 165 456 169
rect 464 165 466 169
rect 480 165 482 169
rect 490 165 492 169
rect 500 165 502 169
rect 516 165 518 169
rect 526 165 528 169
rect 543 165 545 169
rect 553 165 555 169
rect 563 165 565 169
rect 573 165 575 169
rect 589 165 591 169
rect 599 165 601 169
rect 609 165 611 169
rect -332 97 -330 101
rect -322 97 -320 101
rect -305 97 -303 101
rect -295 97 -293 101
rect -285 97 -283 101
rect -275 97 -273 101
rect -259 97 -257 101
rect -249 97 -247 101
rect -239 97 -237 101
rect -223 97 -221 101
rect -213 97 -211 101
rect -196 97 -194 101
rect -186 97 -184 101
rect -176 97 -174 101
rect -166 97 -164 101
rect -150 97 -148 101
rect -140 97 -138 101
rect -130 97 -128 101
rect -114 80 -112 84
rect -101 80 -99 84
rect -83 80 -81 84
rect -73 80 -71 84
rect -54 80 -52 84
rect -34 80 -32 84
rect 35 80 37 84
rect 48 80 50 84
rect 66 80 68 84
rect 76 80 78 84
rect 95 80 97 84
rect 115 80 117 84
rect 184 80 186 84
rect 197 80 199 84
rect 215 80 217 84
rect 225 80 227 84
rect 244 80 246 84
rect 264 80 266 84
rect 333 80 335 84
rect 346 80 348 84
rect 364 80 366 84
rect 374 80 376 84
rect 390 80 392 84
rect 405 80 407 84
rect 561 97 563 101
rect 571 97 573 101
rect 588 97 590 101
rect 598 97 600 101
rect 608 97 610 101
rect 618 97 620 101
rect 634 97 636 101
rect 644 97 646 101
rect 654 97 656 101
rect 465 80 467 84
rect 478 80 480 84
rect 496 80 498 84
rect 506 80 508 84
rect 523 80 525 84
rect 537 80 539 84
rect -10 73 -8 77
rect 0 73 2 77
rect 10 73 12 77
rect 139 73 141 77
rect 149 73 151 77
rect 159 73 161 77
rect 288 73 290 77
rect 298 73 300 77
rect 308 73 310 77
rect 427 73 429 77
rect 437 73 439 77
rect 447 73 449 77
rect -279 -22 -277 -18
rect -269 -22 -267 -18
rect -252 -22 -250 -18
rect -242 -22 -240 -18
rect -232 -22 -230 -18
rect -222 -22 -220 -18
rect -206 -22 -204 -18
rect -196 -22 -194 -18
rect -186 -22 -184 -18
rect 38 -22 40 -18
rect 48 -22 50 -18
rect 58 -22 60 -18
rect 88 -22 90 -18
rect 98 -22 100 -18
rect 108 -22 110 -18
rect 133 -22 135 -18
rect 143 -22 145 -18
rect 153 -22 155 -18
rect 177 -22 179 -18
rect 187 -22 189 -18
rect 197 -22 199 -18
rect 215 -22 217 -18
rect 240 -22 242 -18
rect 250 -22 252 -18
rect 260 -22 262 -18
rect 278 -22 280 -18
rect 305 -22 307 -18
rect 315 -22 317 -18
rect 325 -22 327 -18
rect 336 -22 338 -18
rect 354 -22 356 -18
rect 380 -22 382 -18
rect 390 -22 392 -18
rect 400 -22 402 -18
rect 418 -22 420 -18
rect 434 -22 436 -18
rect 444 -22 446 -18
rect 454 -22 456 -18
rect 479 -22 481 -18
rect 489 -22 491 -18
rect 499 -22 501 -18
rect 510 -22 512 -18
rect 528 -22 530 -18
rect 545 -22 547 -18
rect 555 -22 557 -18
rect 572 -22 574 -18
rect 582 -22 584 -18
rect 592 -22 594 -18
rect 602 -22 604 -18
rect 618 -22 620 -18
rect 628 -22 630 -18
rect 638 -22 640 -18
rect -170 -39 -168 -35
rect -157 -39 -155 -35
rect -139 -39 -137 -35
rect -129 -39 -127 -35
rect -110 -39 -108 -35
rect -90 -39 -88 -35
rect -66 -39 -64 -35
rect -53 -39 -51 -35
rect -35 -39 -33 -35
rect -25 -39 -23 -35
rect -6 -39 -4 -35
rect 14 -39 16 -35
<< ptransistor >>
rect -257 198 -255 206
rect -247 198 -245 206
rect -230 198 -228 206
rect -220 198 -218 206
rect -210 198 -208 206
rect -200 198 -198 206
rect -184 198 -182 206
rect -174 198 -172 206
rect -164 198 -162 206
rect -148 198 -146 206
rect -138 198 -136 206
rect -121 198 -119 206
rect -111 198 -109 206
rect -101 198 -99 206
rect -91 198 -89 206
rect -75 198 -73 206
rect -65 198 -63 206
rect -55 198 -53 206
rect -29 198 -27 206
rect -19 198 -17 206
rect -2 198 0 206
rect 8 198 10 206
rect 18 198 20 206
rect 28 198 30 206
rect 44 198 46 206
rect 54 198 56 206
rect 64 198 66 206
rect 80 198 82 206
rect 90 198 92 206
rect 107 198 109 206
rect 117 198 119 206
rect 127 198 129 206
rect 137 198 139 206
rect 153 198 155 206
rect 163 198 165 206
rect 173 198 175 206
rect 189 198 191 206
rect 199 198 201 206
rect 216 198 218 206
rect 226 198 228 206
rect 236 198 238 206
rect 246 198 248 206
rect 262 198 264 206
rect 272 198 274 206
rect 282 198 284 206
rect 298 198 300 206
rect 308 198 310 206
rect 325 198 327 206
rect 335 198 337 206
rect 345 198 347 206
rect 355 198 357 206
rect 371 198 373 206
rect 381 198 383 206
rect 391 198 393 206
rect 407 198 409 206
rect 417 198 419 206
rect 434 198 436 206
rect 444 198 446 206
rect 454 198 456 206
rect 464 198 466 206
rect 480 198 482 206
rect 490 198 492 206
rect 500 198 502 206
rect 516 198 518 206
rect 526 198 528 206
rect 543 198 545 206
rect 553 198 555 206
rect 563 198 565 206
rect 573 198 575 206
rect 589 198 591 206
rect 599 198 601 206
rect 609 198 611 206
rect -332 130 -330 138
rect -322 130 -320 138
rect -305 130 -303 138
rect -295 130 -293 138
rect -285 130 -283 138
rect -275 130 -273 138
rect -259 130 -257 138
rect -249 130 -247 138
rect -239 130 -237 138
rect -223 130 -221 138
rect -213 130 -211 138
rect -196 130 -194 138
rect -186 130 -184 138
rect -176 130 -174 138
rect -166 130 -164 138
rect -150 130 -148 138
rect -140 130 -138 138
rect -130 130 -128 138
rect -114 130 -112 138
rect -101 130 -99 138
rect -83 130 -81 138
rect -73 130 -71 138
rect -54 130 -52 138
rect -34 130 -32 138
rect -10 130 -8 138
rect 0 130 2 138
rect 10 130 12 138
rect 35 130 37 138
rect 48 130 50 138
rect 66 130 68 138
rect 76 130 78 138
rect 95 130 97 138
rect 115 130 117 138
rect 139 130 141 138
rect 149 130 151 138
rect 159 130 161 138
rect 184 130 186 138
rect 197 130 199 138
rect 215 130 217 138
rect 225 130 227 138
rect 244 130 246 138
rect 264 130 266 138
rect 288 130 290 138
rect 298 130 300 138
rect 308 130 310 138
rect 333 130 335 138
rect 346 130 348 138
rect 364 130 366 138
rect 374 130 376 138
rect 390 130 392 138
rect 405 130 407 138
rect 427 130 429 138
rect 437 130 439 138
rect 447 130 449 138
rect 465 130 467 138
rect 478 130 480 138
rect 496 130 498 138
rect 506 130 508 138
rect 523 130 525 138
rect 537 130 539 138
rect 561 130 563 138
rect 571 130 573 138
rect 588 130 590 138
rect 598 130 600 138
rect 608 130 610 138
rect 618 130 620 138
rect 634 130 636 138
rect 644 130 646 138
rect 654 130 656 138
rect -279 11 -277 19
rect -269 11 -267 19
rect -252 11 -250 19
rect -242 11 -240 19
rect -232 11 -230 19
rect -222 11 -220 19
rect -206 11 -204 19
rect -196 11 -194 19
rect -186 11 -184 19
rect -170 11 -168 19
rect -157 11 -155 19
rect -139 11 -137 19
rect -129 11 -127 19
rect -110 11 -108 19
rect -90 11 -88 19
rect -66 11 -64 19
rect -53 11 -51 19
rect -35 11 -33 19
rect -25 11 -23 19
rect -6 11 -4 19
rect 14 11 16 19
rect 38 11 40 19
rect 48 11 50 19
rect 58 11 60 19
rect 88 11 90 19
rect 98 11 100 19
rect 108 11 110 19
rect 133 11 135 19
rect 143 11 145 19
rect 153 11 155 19
rect 177 11 179 19
rect 187 11 189 19
rect 197 11 199 19
rect 215 11 217 19
rect 240 11 242 19
rect 250 11 252 19
rect 260 11 262 19
rect 278 11 280 19
rect 305 11 307 19
rect 315 11 317 19
rect 325 11 327 19
rect 336 11 338 19
rect 354 11 356 19
rect 380 11 382 19
rect 390 11 392 19
rect 400 11 402 19
rect 418 11 420 19
rect 434 11 436 19
rect 444 11 446 19
rect 454 11 456 19
rect 479 11 481 19
rect 489 11 491 19
rect 499 11 501 19
rect 510 11 512 19
rect 528 11 530 19
rect 545 11 547 19
rect 555 11 557 19
rect 572 11 574 19
rect 582 11 584 19
rect 592 11 594 19
rect 602 11 604 19
rect 618 11 620 19
rect 628 11 630 19
rect 638 11 640 19
<< ndiffusion >>
rect -258 165 -257 169
rect -255 165 -247 169
rect -245 165 -243 169
rect -231 165 -230 169
rect -228 165 -220 169
rect -218 165 -216 169
rect -212 165 -210 169
rect -208 165 -200 169
rect -198 165 -197 169
rect -185 165 -184 169
rect -182 165 -174 169
rect -172 165 -170 169
rect -166 165 -164 169
rect -162 165 -161 169
rect -149 165 -148 169
rect -146 165 -138 169
rect -136 165 -134 169
rect -122 165 -121 169
rect -119 165 -111 169
rect -109 165 -107 169
rect -103 165 -101 169
rect -99 165 -91 169
rect -89 165 -88 169
rect -76 165 -75 169
rect -73 165 -65 169
rect -63 165 -61 169
rect -57 165 -55 169
rect -53 165 -52 169
rect -30 165 -29 169
rect -27 165 -19 169
rect -17 165 -15 169
rect -3 165 -2 169
rect 0 165 8 169
rect 10 165 12 169
rect 16 165 18 169
rect 20 165 28 169
rect 30 165 31 169
rect 43 165 44 169
rect 46 165 54 169
rect 56 165 58 169
rect 62 165 64 169
rect 66 165 67 169
rect 79 165 80 169
rect 82 165 90 169
rect 92 165 94 169
rect 106 165 107 169
rect 109 165 117 169
rect 119 165 121 169
rect 125 165 127 169
rect 129 165 137 169
rect 139 165 140 169
rect 152 165 153 169
rect 155 165 163 169
rect 165 165 167 169
rect 171 165 173 169
rect 175 165 176 169
rect 188 165 189 169
rect 191 165 199 169
rect 201 165 203 169
rect 215 165 216 169
rect 218 165 226 169
rect 228 165 230 169
rect 234 165 236 169
rect 238 165 246 169
rect 248 165 249 169
rect 261 165 262 169
rect 264 165 272 169
rect 274 165 276 169
rect 280 165 282 169
rect 284 165 285 169
rect 297 165 298 169
rect 300 165 308 169
rect 310 165 312 169
rect 324 165 325 169
rect 327 165 335 169
rect 337 165 339 169
rect 343 165 345 169
rect 347 165 355 169
rect 357 165 358 169
rect 370 165 371 169
rect 373 165 381 169
rect 383 165 385 169
rect 389 165 391 169
rect 393 165 394 169
rect 406 165 407 169
rect 409 165 417 169
rect 419 165 421 169
rect 433 165 434 169
rect 436 165 444 169
rect 446 165 448 169
rect 452 165 454 169
rect 456 165 464 169
rect 466 165 467 169
rect 479 165 480 169
rect 482 165 490 169
rect 492 165 494 169
rect 498 165 500 169
rect 502 165 503 169
rect 515 165 516 169
rect 518 165 526 169
rect 528 165 530 169
rect 542 165 543 169
rect 545 165 553 169
rect 555 165 557 169
rect 561 165 563 169
rect 565 165 573 169
rect 575 165 576 169
rect 588 165 589 169
rect 591 165 599 169
rect 601 165 603 169
rect 607 165 609 169
rect 611 165 612 169
rect -333 97 -332 101
rect -330 97 -322 101
rect -320 97 -318 101
rect -306 97 -305 101
rect -303 97 -295 101
rect -293 97 -291 101
rect -287 97 -285 101
rect -283 97 -275 101
rect -273 97 -272 101
rect -260 97 -259 101
rect -257 97 -249 101
rect -247 97 -245 101
rect -241 97 -239 101
rect -237 97 -236 101
rect -224 97 -223 101
rect -221 97 -213 101
rect -211 97 -209 101
rect -197 97 -196 101
rect -194 97 -186 101
rect -184 97 -182 101
rect -178 97 -176 101
rect -174 97 -166 101
rect -164 97 -163 101
rect -151 97 -150 101
rect -148 97 -140 101
rect -138 97 -136 101
rect -132 97 -130 101
rect -128 97 -127 101
rect -115 80 -114 84
rect -112 80 -109 84
rect -105 80 -101 84
rect -99 80 -98 84
rect -84 80 -83 84
rect -81 80 -79 84
rect -75 80 -73 84
rect -71 80 -69 84
rect -65 80 -54 84
rect -52 80 -50 84
rect -46 80 -34 84
rect -32 80 -31 84
rect 34 80 35 84
rect 37 80 40 84
rect 44 80 48 84
rect 50 80 51 84
rect 65 80 66 84
rect 68 80 70 84
rect 74 80 76 84
rect 78 80 80 84
rect 84 80 95 84
rect 97 80 99 84
rect 103 80 115 84
rect 117 80 118 84
rect 183 80 184 84
rect 186 80 189 84
rect 193 80 197 84
rect 199 80 200 84
rect 214 80 215 84
rect 217 80 219 84
rect 223 80 225 84
rect 227 80 229 84
rect 233 80 244 84
rect 246 80 248 84
rect 252 80 264 84
rect 266 80 267 84
rect 332 80 333 84
rect 335 80 338 84
rect 342 80 346 84
rect 348 80 349 84
rect 363 80 364 84
rect 366 80 368 84
rect 372 80 374 84
rect 376 80 378 84
rect 382 80 390 84
rect 392 80 394 84
rect 398 80 405 84
rect 407 80 408 84
rect 560 97 561 101
rect 563 97 571 101
rect 573 97 575 101
rect 587 97 588 101
rect 590 97 598 101
rect 600 97 602 101
rect 606 97 608 101
rect 610 97 618 101
rect 620 97 621 101
rect 633 97 634 101
rect 636 97 644 101
rect 646 97 648 101
rect 652 97 654 101
rect 656 97 657 101
rect 464 80 465 84
rect 467 80 470 84
rect 474 80 478 84
rect 480 80 481 84
rect 495 80 496 84
rect 498 80 500 84
rect 504 80 506 84
rect 508 80 510 84
rect 514 80 523 84
rect 525 80 527 84
rect 531 80 537 84
rect 539 80 540 84
rect -11 73 -10 77
rect -8 73 0 77
rect 2 73 4 77
rect 8 73 10 77
rect 12 73 13 77
rect 138 73 139 77
rect 141 73 149 77
rect 151 73 153 77
rect 157 73 159 77
rect 161 73 162 77
rect 287 73 288 77
rect 290 73 298 77
rect 300 73 302 77
rect 306 73 308 77
rect 310 73 311 77
rect 426 73 427 77
rect 429 73 437 77
rect 439 73 441 77
rect 445 73 447 77
rect 449 73 450 77
rect -280 -22 -279 -18
rect -277 -22 -269 -18
rect -267 -22 -265 -18
rect -253 -22 -252 -18
rect -250 -22 -242 -18
rect -240 -22 -238 -18
rect -234 -22 -232 -18
rect -230 -22 -222 -18
rect -220 -22 -219 -18
rect -207 -22 -206 -18
rect -204 -22 -196 -18
rect -194 -22 -192 -18
rect -188 -22 -186 -18
rect -184 -22 -183 -18
rect 37 -22 38 -18
rect 40 -22 48 -18
rect 50 -22 52 -18
rect 56 -22 58 -18
rect 60 -22 61 -18
rect 87 -22 88 -18
rect 90 -22 92 -18
rect 96 -22 98 -18
rect 100 -22 102 -18
rect 106 -22 108 -18
rect 110 -22 111 -18
rect 132 -22 133 -18
rect 135 -22 143 -18
rect 145 -22 147 -18
rect 151 -22 153 -18
rect 155 -22 156 -18
rect 176 -22 177 -18
rect 179 -22 187 -18
rect 189 -22 197 -18
rect 199 -22 200 -18
rect 209 -22 210 -18
rect 214 -22 215 -18
rect 217 -22 218 -18
rect 239 -22 240 -18
rect 242 -22 244 -18
rect 248 -22 250 -18
rect 252 -22 254 -18
rect 258 -22 260 -18
rect 262 -22 263 -18
rect 272 -22 273 -18
rect 277 -22 278 -18
rect 280 -22 281 -18
rect 304 -22 305 -18
rect 307 -22 315 -18
rect 317 -22 325 -18
rect 327 -22 336 -18
rect 338 -22 339 -18
rect 348 -22 349 -18
rect 353 -22 354 -18
rect 356 -22 357 -18
rect 379 -22 380 -18
rect 382 -22 390 -18
rect 392 -22 400 -18
rect 402 -22 403 -18
rect 412 -22 413 -18
rect 417 -22 418 -18
rect 420 -22 421 -18
rect 433 -22 434 -18
rect 436 -22 444 -18
rect 446 -22 448 -18
rect 452 -22 454 -18
rect 456 -22 457 -18
rect 478 -22 479 -18
rect 481 -22 483 -18
rect 487 -22 489 -18
rect 491 -22 493 -18
rect 497 -22 499 -18
rect 501 -22 504 -18
rect 508 -22 510 -18
rect 512 -22 513 -18
rect 522 -22 523 -18
rect 527 -22 528 -18
rect 530 -22 531 -18
rect 544 -22 545 -18
rect 547 -22 555 -18
rect 557 -22 559 -18
rect 571 -22 572 -18
rect 574 -22 582 -18
rect 584 -22 586 -18
rect 590 -22 592 -18
rect 594 -22 602 -18
rect 604 -22 605 -18
rect 617 -22 618 -18
rect 620 -22 628 -18
rect 630 -22 632 -18
rect 636 -22 638 -18
rect 640 -22 641 -18
rect -171 -39 -170 -35
rect -168 -39 -165 -35
rect -161 -39 -157 -35
rect -155 -39 -154 -35
rect -140 -39 -139 -35
rect -137 -39 -135 -35
rect -131 -39 -129 -35
rect -127 -39 -125 -35
rect -121 -39 -110 -35
rect -108 -39 -106 -35
rect -102 -39 -90 -35
rect -88 -39 -87 -35
rect -67 -39 -66 -35
rect -64 -39 -61 -35
rect -57 -39 -53 -35
rect -51 -39 -50 -35
rect -36 -39 -35 -35
rect -33 -39 -31 -35
rect -27 -39 -25 -35
rect -23 -39 -21 -35
rect -17 -39 -6 -35
rect -4 -39 -2 -35
rect 2 -39 14 -35
rect 16 -39 17 -35
<< pdiffusion >>
rect -258 198 -257 206
rect -255 198 -253 206
rect -249 198 -247 206
rect -245 198 -240 206
rect -236 198 -230 206
rect -228 198 -226 206
rect -222 198 -220 206
rect -218 198 -216 206
rect -212 198 -210 206
rect -208 198 -206 206
rect -202 198 -200 206
rect -198 198 -193 206
rect -189 198 -184 206
rect -182 198 -180 206
rect -176 198 -174 206
rect -172 198 -170 206
rect -166 198 -164 206
rect -162 198 -161 206
rect -149 198 -148 206
rect -146 198 -144 206
rect -140 198 -138 206
rect -136 198 -131 206
rect -127 198 -121 206
rect -119 198 -117 206
rect -113 198 -111 206
rect -109 198 -107 206
rect -103 198 -101 206
rect -99 198 -97 206
rect -93 198 -91 206
rect -89 198 -84 206
rect -80 198 -75 206
rect -73 198 -71 206
rect -67 198 -65 206
rect -63 198 -61 206
rect -57 198 -55 206
rect -53 198 -52 206
rect -30 198 -29 206
rect -27 198 -25 206
rect -21 198 -19 206
rect -17 198 -12 206
rect -8 198 -2 206
rect 0 198 2 206
rect 6 198 8 206
rect 10 198 12 206
rect 16 198 18 206
rect 20 198 22 206
rect 26 198 28 206
rect 30 198 35 206
rect 39 198 44 206
rect 46 198 48 206
rect 52 198 54 206
rect 56 198 58 206
rect 62 198 64 206
rect 66 198 67 206
rect 79 198 80 206
rect 82 198 84 206
rect 88 198 90 206
rect 92 198 97 206
rect 101 198 107 206
rect 109 198 111 206
rect 115 198 117 206
rect 119 198 121 206
rect 125 198 127 206
rect 129 198 131 206
rect 135 198 137 206
rect 139 198 144 206
rect 148 198 153 206
rect 155 198 157 206
rect 161 198 163 206
rect 165 198 167 206
rect 171 198 173 206
rect 175 198 176 206
rect 188 198 189 206
rect 191 198 193 206
rect 197 198 199 206
rect 201 198 206 206
rect 210 198 216 206
rect 218 198 220 206
rect 224 198 226 206
rect 228 198 230 206
rect 234 198 236 206
rect 238 198 240 206
rect 244 198 246 206
rect 248 198 253 206
rect 257 198 262 206
rect 264 198 266 206
rect 270 198 272 206
rect 274 198 276 206
rect 280 198 282 206
rect 284 198 285 206
rect 297 198 298 206
rect 300 198 302 206
rect 306 198 308 206
rect 310 198 315 206
rect 319 198 325 206
rect 327 198 329 206
rect 333 198 335 206
rect 337 198 339 206
rect 343 198 345 206
rect 347 198 349 206
rect 353 198 355 206
rect 357 198 362 206
rect 366 198 371 206
rect 373 198 375 206
rect 379 198 381 206
rect 383 198 385 206
rect 389 198 391 206
rect 393 198 394 206
rect 406 198 407 206
rect 409 198 411 206
rect 415 198 417 206
rect 419 198 424 206
rect 428 198 434 206
rect 436 198 438 206
rect 442 198 444 206
rect 446 198 448 206
rect 452 198 454 206
rect 456 198 458 206
rect 462 198 464 206
rect 466 198 471 206
rect 475 198 480 206
rect 482 198 484 206
rect 488 198 490 206
rect 492 198 494 206
rect 498 198 500 206
rect 502 198 503 206
rect 515 198 516 206
rect 518 198 520 206
rect 524 198 526 206
rect 528 198 533 206
rect 537 198 543 206
rect 545 198 547 206
rect 551 198 553 206
rect 555 198 557 206
rect 561 198 563 206
rect 565 198 567 206
rect 571 198 573 206
rect 575 198 580 206
rect 584 198 589 206
rect 591 198 593 206
rect 597 198 599 206
rect 601 198 603 206
rect 607 198 609 206
rect 611 198 612 206
rect -333 130 -332 138
rect -330 130 -328 138
rect -324 130 -322 138
rect -320 130 -315 138
rect -311 130 -305 138
rect -303 130 -301 138
rect -297 130 -295 138
rect -293 130 -291 138
rect -287 130 -285 138
rect -283 130 -281 138
rect -277 130 -275 138
rect -273 130 -268 138
rect -264 130 -259 138
rect -257 130 -255 138
rect -251 130 -249 138
rect -247 130 -245 138
rect -241 130 -239 138
rect -237 130 -236 138
rect -224 130 -223 138
rect -221 130 -219 138
rect -215 130 -213 138
rect -211 130 -206 138
rect -202 130 -196 138
rect -194 130 -192 138
rect -188 130 -186 138
rect -184 130 -182 138
rect -178 130 -176 138
rect -174 130 -172 138
rect -168 130 -166 138
rect -164 130 -159 138
rect -155 130 -150 138
rect -148 130 -146 138
rect -142 130 -140 138
rect -138 130 -136 138
rect -132 130 -130 138
rect -128 130 -127 138
rect -115 130 -114 138
rect -112 130 -106 138
rect -102 130 -101 138
rect -99 130 -98 138
rect -84 130 -83 138
rect -81 130 -73 138
rect -71 130 -69 138
rect -65 130 -54 138
rect -52 130 -34 138
rect -32 130 -31 138
rect -11 130 -10 138
rect -8 130 -6 138
rect -2 130 0 138
rect 2 130 4 138
rect 8 130 10 138
rect 12 130 13 138
rect 34 130 35 138
rect 37 130 43 138
rect 47 130 48 138
rect 50 130 51 138
rect 65 130 66 138
rect 68 130 76 138
rect 78 130 80 138
rect 84 130 95 138
rect 97 130 115 138
rect 117 130 118 138
rect 138 130 139 138
rect 141 130 143 138
rect 147 130 149 138
rect 151 130 153 138
rect 157 130 159 138
rect 161 130 162 138
rect 183 130 184 138
rect 186 130 192 138
rect 196 130 197 138
rect 199 130 200 138
rect 214 130 215 138
rect 217 130 225 138
rect 227 130 229 138
rect 233 130 244 138
rect 246 130 264 138
rect 266 130 267 138
rect 287 130 288 138
rect 290 130 292 138
rect 296 130 298 138
rect 300 130 302 138
rect 306 130 308 138
rect 310 130 311 138
rect 332 130 333 138
rect 335 130 341 138
rect 345 130 346 138
rect 348 130 349 138
rect 363 130 364 138
rect 366 130 374 138
rect 376 130 378 138
rect 382 130 390 138
rect 392 130 405 138
rect 407 130 408 138
rect 426 130 427 138
rect 429 130 431 138
rect 435 130 437 138
rect 439 130 441 138
rect 445 130 447 138
rect 449 130 450 138
rect 464 130 465 138
rect 467 130 473 138
rect 477 130 478 138
rect 480 130 481 138
rect 495 130 496 138
rect 498 130 506 138
rect 508 130 510 138
rect 514 130 523 138
rect 525 130 537 138
rect 539 130 540 138
rect 560 130 561 138
rect 563 130 565 138
rect 569 130 571 138
rect 573 130 578 138
rect 582 130 588 138
rect 590 130 592 138
rect 596 130 598 138
rect 600 130 602 138
rect 606 130 608 138
rect 610 130 612 138
rect 616 130 618 138
rect 620 130 625 138
rect 629 130 634 138
rect 636 130 638 138
rect 642 130 644 138
rect 646 130 648 138
rect 652 130 654 138
rect 656 130 657 138
rect -280 11 -279 19
rect -277 11 -275 19
rect -271 11 -269 19
rect -267 11 -262 19
rect -258 11 -252 19
rect -250 11 -248 19
rect -244 11 -242 19
rect -240 11 -238 19
rect -234 11 -232 19
rect -230 11 -228 19
rect -224 11 -222 19
rect -220 11 -215 19
rect -211 11 -206 19
rect -204 11 -202 19
rect -198 11 -196 19
rect -194 11 -192 19
rect -188 11 -186 19
rect -184 11 -183 19
rect -171 11 -170 19
rect -168 11 -162 19
rect -158 11 -157 19
rect -155 11 -154 19
rect -140 11 -139 19
rect -137 11 -129 19
rect -127 11 -125 19
rect -121 11 -110 19
rect -108 11 -90 19
rect -88 11 -87 19
rect -67 11 -66 19
rect -64 11 -58 19
rect -54 11 -53 19
rect -51 11 -50 19
rect -36 11 -35 19
rect -33 11 -25 19
rect -23 11 -21 19
rect -17 11 -6 19
rect -4 11 14 19
rect 16 11 17 19
rect 37 11 38 19
rect 40 11 42 19
rect 46 11 48 19
rect 50 11 52 19
rect 56 11 58 19
rect 60 11 61 19
rect 87 11 88 19
rect 90 11 98 19
rect 100 11 102 19
rect 106 11 108 19
rect 110 11 111 19
rect 132 11 133 19
rect 135 11 137 19
rect 141 11 143 19
rect 145 11 147 19
rect 151 11 153 19
rect 155 11 156 19
rect 176 11 177 19
rect 179 11 181 19
rect 185 11 187 19
rect 189 11 191 19
rect 195 11 197 19
rect 199 11 200 19
rect 208 11 210 19
rect 214 11 215 19
rect 217 11 218 19
rect 239 11 240 19
rect 242 11 250 19
rect 252 11 260 19
rect 262 11 263 19
rect 272 11 273 19
rect 277 11 278 19
rect 280 11 281 19
rect 304 11 305 19
rect 307 11 309 19
rect 313 11 315 19
rect 317 11 319 19
rect 323 11 325 19
rect 327 11 329 19
rect 333 11 336 19
rect 338 11 339 19
rect 348 11 349 19
rect 353 11 354 19
rect 356 11 357 19
rect 379 11 380 19
rect 382 11 384 19
rect 388 11 390 19
rect 392 11 394 19
rect 398 11 400 19
rect 402 11 403 19
rect 411 11 413 19
rect 417 11 418 19
rect 420 11 421 19
rect 433 11 434 19
rect 436 11 438 19
rect 442 11 444 19
rect 446 11 448 19
rect 452 11 454 19
rect 456 11 457 19
rect 478 11 479 19
rect 481 11 489 19
rect 491 11 499 19
rect 501 11 510 19
rect 512 11 513 19
rect 522 11 523 19
rect 527 11 528 19
rect 530 11 531 19
rect 544 11 545 19
rect 547 11 549 19
rect 553 11 555 19
rect 557 11 562 19
rect 566 11 572 19
rect 574 11 576 19
rect 580 11 582 19
rect 584 11 586 19
rect 590 11 592 19
rect 594 11 596 19
rect 600 11 602 19
rect 604 11 609 19
rect 613 11 618 19
rect 620 11 622 19
rect 626 11 628 19
rect 630 11 632 19
rect 636 11 638 19
rect 640 11 641 19
<< ndcontact >>
rect -262 165 -258 169
rect -243 165 -239 169
rect -235 165 -231 169
rect -216 165 -212 169
rect -197 165 -193 169
rect -189 165 -185 169
rect -170 165 -166 169
rect -161 165 -157 169
rect -153 165 -149 169
rect -134 165 -130 169
rect -126 165 -122 169
rect -107 165 -103 169
rect -88 165 -84 169
rect -80 165 -76 169
rect -61 165 -57 169
rect -52 165 -48 169
rect -34 165 -30 169
rect -15 165 -11 169
rect -7 165 -3 169
rect 12 165 16 169
rect 31 165 35 169
rect 39 165 43 169
rect 58 165 62 169
rect 67 165 71 169
rect 75 165 79 169
rect 94 165 98 169
rect 102 165 106 169
rect 121 165 125 169
rect 140 165 144 169
rect 148 165 152 169
rect 167 165 171 169
rect 176 165 180 169
rect 184 165 188 169
rect 203 165 207 169
rect 211 165 215 169
rect 230 165 234 169
rect 249 165 253 169
rect 257 165 261 169
rect 276 165 280 169
rect 285 165 289 169
rect 293 165 297 169
rect 312 165 316 169
rect 320 165 324 169
rect 339 165 343 169
rect 358 165 362 169
rect 366 165 370 169
rect 385 165 389 169
rect 394 165 398 169
rect 402 165 406 169
rect 421 165 425 169
rect 429 165 433 169
rect 448 165 452 169
rect 467 165 471 169
rect 475 165 479 169
rect 494 165 498 169
rect 503 165 507 169
rect 511 165 515 169
rect 530 165 534 169
rect 538 165 542 169
rect 557 165 561 169
rect 576 165 580 169
rect 584 165 588 169
rect 603 165 607 169
rect 612 165 616 169
rect -337 97 -333 101
rect -318 97 -314 101
rect -310 97 -306 101
rect -291 97 -287 101
rect -272 97 -268 101
rect -264 97 -260 101
rect -245 97 -241 101
rect -236 97 -232 101
rect -228 97 -224 101
rect -209 97 -205 101
rect -201 97 -197 101
rect -182 97 -178 101
rect -163 97 -159 101
rect -155 97 -151 101
rect -136 97 -132 101
rect -127 97 -123 101
rect -119 80 -115 84
rect -109 80 -105 84
rect -98 80 -94 84
rect -88 80 -84 84
rect -79 80 -75 84
rect -69 80 -65 84
rect -50 80 -46 84
rect -31 80 -27 84
rect 30 80 34 84
rect 40 80 44 84
rect 51 80 55 84
rect 61 80 65 84
rect 70 80 74 84
rect 80 80 84 84
rect 99 80 103 84
rect 118 80 122 84
rect 179 80 183 84
rect 189 80 193 84
rect 200 80 204 84
rect 210 80 214 84
rect 219 80 223 84
rect 229 80 233 84
rect 248 80 252 84
rect 267 80 271 84
rect 328 80 332 84
rect 338 80 342 84
rect 349 80 353 84
rect 359 80 363 84
rect 368 80 372 84
rect 378 80 382 84
rect 394 80 398 84
rect 408 80 412 84
rect 556 97 560 101
rect 575 97 579 101
rect 583 97 587 101
rect 602 97 606 101
rect 621 97 625 101
rect 629 97 633 101
rect 648 97 652 101
rect 657 97 661 101
rect 460 80 464 84
rect 470 80 474 84
rect 481 80 485 84
rect 491 80 495 84
rect 500 80 504 84
rect 510 80 514 84
rect 527 80 531 84
rect 540 80 544 84
rect -15 73 -11 77
rect 4 73 8 77
rect 13 73 17 77
rect 134 73 138 77
rect 153 73 157 77
rect 162 73 166 77
rect 283 73 287 77
rect 302 73 306 77
rect 311 73 315 77
rect 422 73 426 77
rect 441 73 445 77
rect 450 73 454 77
rect -284 -22 -280 -18
rect -265 -22 -261 -18
rect -257 -22 -253 -18
rect -238 -22 -234 -18
rect -219 -22 -215 -18
rect -211 -22 -207 -18
rect -192 -22 -188 -18
rect -183 -22 -179 -18
rect 33 -22 37 -18
rect 52 -22 56 -18
rect 61 -22 65 -18
rect 83 -22 87 -18
rect 92 -22 96 -18
rect 102 -22 106 -18
rect 111 -22 115 -18
rect 128 -22 132 -18
rect 147 -22 151 -18
rect 156 -22 160 -18
rect 172 -22 176 -18
rect 200 -22 204 -18
rect 210 -22 214 -18
rect 218 -22 222 -18
rect 235 -22 239 -18
rect 244 -22 248 -18
rect 254 -22 258 -18
rect 263 -22 267 -18
rect 273 -22 277 -18
rect 281 -22 285 -18
rect 300 -22 304 -18
rect 339 -22 343 -18
rect 349 -22 353 -18
rect 357 -22 361 -18
rect 375 -22 379 -18
rect 403 -22 407 -18
rect 413 -22 417 -18
rect 421 -22 425 -18
rect 429 -22 433 -18
rect 448 -22 452 -18
rect 457 -22 461 -18
rect 474 -22 478 -18
rect 483 -22 487 -18
rect 493 -22 497 -18
rect 504 -22 508 -18
rect 513 -22 517 -18
rect 523 -22 527 -18
rect 531 -22 535 -18
rect 540 -22 544 -18
rect 559 -22 563 -18
rect 567 -22 571 -18
rect 586 -22 590 -18
rect 605 -22 609 -18
rect 613 -22 617 -18
rect 632 -22 636 -18
rect 641 -22 645 -18
rect -175 -39 -171 -35
rect -165 -39 -161 -35
rect -154 -39 -150 -35
rect -144 -39 -140 -35
rect -135 -39 -131 -35
rect -125 -39 -121 -35
rect -106 -39 -102 -35
rect -87 -39 -83 -35
rect -71 -39 -67 -35
rect -61 -39 -57 -35
rect -50 -39 -46 -35
rect -40 -39 -36 -35
rect -31 -39 -27 -35
rect -21 -39 -17 -35
rect -2 -39 2 -35
rect 17 -39 21 -35
<< pdcontact >>
rect -262 198 -258 206
rect -253 198 -249 206
rect -240 198 -236 206
rect -226 198 -222 206
rect -216 198 -212 206
rect -206 198 -202 206
rect -193 198 -189 206
rect -180 198 -176 206
rect -170 198 -166 206
rect -161 198 -157 206
rect -153 198 -149 206
rect -144 198 -140 206
rect -131 198 -127 206
rect -117 198 -113 206
rect -107 198 -103 206
rect -97 198 -93 206
rect -84 198 -80 206
rect -71 198 -67 206
rect -61 198 -57 206
rect -52 198 -48 206
rect -34 198 -30 206
rect -25 198 -21 206
rect -12 198 -8 206
rect 2 198 6 206
rect 12 198 16 206
rect 22 198 26 206
rect 35 198 39 206
rect 48 198 52 206
rect 58 198 62 206
rect 67 198 71 206
rect 75 198 79 206
rect 84 198 88 206
rect 97 198 101 206
rect 111 198 115 206
rect 121 198 125 206
rect 131 198 135 206
rect 144 198 148 206
rect 157 198 161 206
rect 167 198 171 206
rect 176 198 180 206
rect 184 198 188 206
rect 193 198 197 206
rect 206 198 210 206
rect 220 198 224 206
rect 230 198 234 206
rect 240 198 244 206
rect 253 198 257 206
rect 266 198 270 206
rect 276 198 280 206
rect 285 198 289 206
rect 293 198 297 206
rect 302 198 306 206
rect 315 198 319 206
rect 329 198 333 206
rect 339 198 343 206
rect 349 198 353 206
rect 362 198 366 206
rect 375 198 379 206
rect 385 198 389 206
rect 394 198 398 206
rect 402 198 406 206
rect 411 198 415 206
rect 424 198 428 206
rect 438 198 442 206
rect 448 198 452 206
rect 458 198 462 206
rect 471 198 475 206
rect 484 198 488 206
rect 494 198 498 206
rect 503 198 507 206
rect 511 198 515 206
rect 520 198 524 206
rect 533 198 537 206
rect 547 198 551 206
rect 557 198 561 206
rect 567 198 571 206
rect 580 198 584 206
rect 593 198 597 206
rect 603 198 607 206
rect 612 198 616 206
rect -337 130 -333 138
rect -328 130 -324 138
rect -315 130 -311 138
rect -301 130 -297 138
rect -291 130 -287 138
rect -281 130 -277 138
rect -268 130 -264 138
rect -255 130 -251 138
rect -245 130 -241 138
rect -236 130 -232 138
rect -228 130 -224 138
rect -219 130 -215 138
rect -206 130 -202 138
rect -192 130 -188 138
rect -182 130 -178 138
rect -172 130 -168 138
rect -159 130 -155 138
rect -146 130 -142 138
rect -136 130 -132 138
rect -127 130 -123 138
rect -119 130 -115 138
rect -106 130 -102 138
rect -98 130 -94 138
rect -88 130 -84 138
rect -69 130 -65 138
rect -31 130 -27 138
rect -15 130 -11 138
rect -6 130 -2 138
rect 4 130 8 138
rect 13 130 17 138
rect 30 130 34 138
rect 43 130 47 138
rect 51 130 55 138
rect 61 130 65 138
rect 80 130 84 138
rect 118 130 122 138
rect 134 130 138 138
rect 143 130 147 138
rect 153 130 157 138
rect 162 130 166 138
rect 179 130 183 138
rect 192 130 196 138
rect 200 130 204 138
rect 210 130 214 138
rect 229 130 233 138
rect 267 130 271 138
rect 283 130 287 138
rect 292 130 296 138
rect 302 130 306 138
rect 311 130 315 138
rect 328 130 332 138
rect 341 130 345 138
rect 349 130 353 138
rect 359 130 363 138
rect 378 130 382 138
rect 408 130 412 138
rect 422 130 426 138
rect 431 130 435 138
rect 441 130 445 138
rect 450 130 454 138
rect 460 130 464 138
rect 473 130 477 138
rect 481 130 485 138
rect 491 130 495 138
rect 510 130 514 138
rect 540 130 544 138
rect 556 130 560 138
rect 565 130 569 138
rect 578 130 582 138
rect 592 130 596 138
rect 602 130 606 138
rect 612 130 616 138
rect 625 130 629 138
rect 638 130 642 138
rect 648 130 652 138
rect 657 130 661 138
rect -284 11 -280 19
rect -275 11 -271 19
rect -262 11 -258 19
rect -248 11 -244 19
rect -238 11 -234 19
rect -228 11 -224 19
rect -215 11 -211 19
rect -202 11 -198 19
rect -192 11 -188 19
rect -183 11 -179 19
rect -175 11 -171 19
rect -162 11 -158 19
rect -154 11 -150 19
rect -144 11 -140 19
rect -125 11 -121 19
rect -87 11 -83 19
rect -71 11 -67 19
rect -58 11 -54 19
rect -50 11 -46 19
rect -40 11 -36 19
rect -21 11 -17 19
rect 17 11 21 19
rect 33 11 37 19
rect 42 11 46 19
rect 52 11 56 19
rect 61 11 65 19
rect 83 11 87 19
rect 102 11 106 19
rect 111 11 115 19
rect 128 11 132 19
rect 137 11 141 19
rect 147 11 151 19
rect 156 11 160 19
rect 172 11 176 19
rect 181 11 185 19
rect 191 11 195 19
rect 200 11 204 19
rect 210 11 214 19
rect 218 11 222 19
rect 235 11 239 19
rect 263 11 267 19
rect 273 11 277 19
rect 281 11 285 19
rect 300 11 304 19
rect 309 11 313 19
rect 319 11 323 19
rect 329 11 333 19
rect 339 11 343 19
rect 349 11 353 19
rect 357 11 361 19
rect 375 11 379 19
rect 384 11 388 19
rect 394 11 398 19
rect 403 11 407 19
rect 413 11 417 19
rect 421 11 425 19
rect 429 11 433 19
rect 438 11 442 19
rect 448 11 452 19
rect 457 11 461 19
rect 474 11 478 19
rect 513 11 517 19
rect 523 11 527 19
rect 531 11 535 19
rect 540 11 544 19
rect 549 11 553 19
rect 562 11 566 19
rect 576 11 580 19
rect 586 11 590 19
rect 596 11 600 19
rect 609 11 613 19
rect 622 11 626 19
rect 632 11 636 19
rect 641 11 645 19
<< psubstratepcontact >>
rect -263 157 -259 161
rect -236 157 -232 161
rect -216 157 -212 161
rect -198 157 -194 161
rect -190 157 -186 161
rect -170 157 -166 161
rect -154 157 -150 161
rect -127 157 -123 161
rect -107 157 -103 161
rect -89 157 -85 161
rect -81 157 -77 161
rect -61 157 -57 161
rect -35 157 -31 161
rect -8 157 -4 161
rect 12 157 16 161
rect 30 157 34 161
rect 38 157 42 161
rect 58 157 62 161
rect 74 157 78 161
rect 101 157 105 161
rect 121 157 125 161
rect 139 157 143 161
rect 147 157 151 161
rect 167 157 171 161
rect 183 157 187 161
rect 210 157 214 161
rect 230 157 234 161
rect 248 157 252 161
rect 256 157 260 161
rect 276 157 280 161
rect 292 157 296 161
rect 319 157 323 161
rect 339 157 343 161
rect 357 157 361 161
rect 365 157 369 161
rect 385 157 389 161
rect 401 157 405 161
rect 428 157 432 161
rect 448 157 452 161
rect 466 157 470 161
rect 474 157 478 161
rect 494 157 498 161
rect 510 157 514 161
rect 537 157 541 161
rect 557 157 561 161
rect 575 157 579 161
rect 583 157 587 161
rect 603 157 607 161
rect -338 89 -334 93
rect -311 89 -307 93
rect -291 89 -287 93
rect -273 89 -269 93
rect -265 89 -261 93
rect -245 89 -241 93
rect -229 89 -225 93
rect -202 89 -198 93
rect -182 89 -178 93
rect -164 89 -160 93
rect -156 89 -152 93
rect -136 89 -132 93
rect 555 89 559 93
rect 582 89 586 93
rect 602 89 606 93
rect 620 89 624 93
rect 628 89 632 93
rect 648 89 652 93
rect -125 65 -121 69
rect -107 65 -103 69
rect -89 65 -85 69
rect -56 65 -52 69
rect -26 65 -22 69
rect -16 65 -12 69
rect 13 65 17 69
rect 24 65 28 69
rect 42 65 46 69
rect 60 65 64 69
rect 93 65 97 69
rect 123 65 127 69
rect 133 65 137 69
rect 162 65 166 69
rect 173 65 177 69
rect 191 65 195 69
rect 209 65 213 69
rect 242 65 246 69
rect 272 65 276 69
rect 282 65 286 69
rect 311 65 315 69
rect 322 65 326 69
rect 340 65 344 69
rect 358 65 362 69
rect 388 65 392 69
rect 413 65 417 69
rect 421 65 425 69
rect 450 65 454 69
rect 458 65 462 69
rect 472 65 476 69
rect 490 65 494 69
rect 523 65 527 69
rect 555 65 559 69
rect -285 -30 -281 -26
rect -258 -30 -254 -26
rect -238 -30 -234 -26
rect -220 -30 -216 -26
rect -212 -30 -208 -26
rect -192 -30 -188 -26
rect 32 -30 36 -26
rect 61 -30 65 -26
rect 82 -30 86 -26
rect 111 -30 115 -26
rect 127 -30 131 -26
rect 156 -30 160 -26
rect 171 -30 175 -26
rect 200 -30 204 -26
rect 222 -30 226 -26
rect 235 -30 239 -26
rect 263 -30 267 -26
rect 285 -30 289 -26
rect 300 -30 304 -26
rect 330 -30 334 -26
rect 361 -30 365 -26
rect 374 -30 378 -26
rect 403 -30 407 -26
rect 425 -30 429 -26
rect 433 -30 437 -26
rect 457 -30 461 -26
rect 474 -30 478 -26
rect 504 -30 508 -26
rect 535 -30 543 -26
rect 566 -30 570 -26
rect 586 -30 590 -26
rect 604 -30 608 -26
rect 612 -30 616 -26
rect 632 -30 636 -26
rect -192 -54 -188 -50
rect -163 -54 -159 -50
rect -145 -54 -141 -50
rect -112 -54 -108 -50
rect -82 -54 -78 -50
rect -61 -54 -57 -50
rect -41 -54 -37 -50
rect -8 -54 -4 -50
rect 22 -54 26 -50
<< nsubstratencontact >>
rect -262 211 -258 215
rect -243 211 -239 215
rect -216 211 -212 215
rect -170 211 -166 215
rect -153 211 -149 215
rect -134 211 -130 215
rect -107 211 -103 215
rect -61 211 -57 215
rect -34 211 -30 215
rect -15 211 -11 215
rect 12 211 16 215
rect 58 211 62 215
rect 75 211 79 215
rect 94 211 98 215
rect 121 211 125 215
rect 167 211 171 215
rect 184 211 188 215
rect 203 211 207 215
rect 230 211 234 215
rect 276 211 280 215
rect 293 211 297 215
rect 312 211 316 215
rect 339 211 343 215
rect 385 211 389 215
rect 402 211 406 215
rect 421 211 425 215
rect 448 211 452 215
rect 494 211 498 215
rect 511 211 515 215
rect 530 211 534 215
rect 557 211 561 215
rect 603 211 607 215
rect -337 143 -333 147
rect -318 143 -314 147
rect -291 143 -287 147
rect -245 143 -241 147
rect -228 143 -224 147
rect -209 143 -205 147
rect -182 143 -178 147
rect -136 143 -132 147
rect -121 143 -117 147
rect -96 143 -92 147
rect -88 143 -84 147
rect -69 143 -65 147
rect -28 143 -24 147
rect -15 143 -11 147
rect 14 143 18 147
rect 28 143 32 147
rect 53 143 57 147
rect 61 143 65 147
rect 80 143 84 147
rect 121 143 125 147
rect 134 143 138 147
rect 163 143 167 147
rect 177 143 181 147
rect 202 143 206 147
rect 210 143 214 147
rect 229 143 233 147
rect 270 143 274 147
rect 283 143 287 147
rect 312 143 316 147
rect 326 143 330 147
rect 351 143 355 147
rect 359 143 363 147
rect 378 143 382 147
rect 411 143 415 147
rect 422 143 426 147
rect 451 143 455 147
rect 467 143 471 147
rect 483 143 487 147
rect 491 143 495 147
rect 510 143 514 147
rect 543 143 547 147
rect 556 143 560 147
rect 575 143 579 147
rect 602 143 606 147
rect 648 143 652 147
rect -284 24 -280 28
rect -265 24 -261 28
rect -238 24 -234 28
rect -192 24 -188 28
rect -177 24 -173 28
rect -152 24 -148 28
rect -144 24 -140 28
rect -125 24 -121 28
rect -84 24 -80 28
rect -73 24 -69 28
rect -48 24 -44 28
rect -40 24 -36 28
rect -21 24 -17 28
rect 20 24 24 28
rect 33 24 37 28
rect 62 24 66 28
rect 83 24 87 28
rect 112 24 116 28
rect 128 24 132 28
rect 157 24 161 28
rect 172 24 176 28
rect 201 24 205 28
rect 220 24 224 28
rect 235 24 239 28
rect 264 24 268 28
rect 283 24 287 28
rect 300 24 304 28
rect 331 24 335 28
rect 359 24 363 28
rect 375 24 379 28
rect 404 24 408 28
rect 429 24 433 28
rect 458 24 462 28
rect 474 24 478 28
rect 505 24 509 28
rect 540 24 544 28
rect 559 24 563 28
rect 586 24 590 28
rect 632 24 636 28
<< polysilicon >>
rect -257 206 -255 222
rect -247 206 -245 209
rect -230 206 -228 209
rect -220 206 -218 209
rect -210 206 -208 209
rect -200 206 -198 209
rect -184 206 -182 209
rect -174 206 -172 209
rect -164 206 -162 222
rect -148 206 -146 222
rect -138 206 -136 209
rect -121 206 -119 209
rect -111 206 -109 209
rect -101 206 -99 209
rect -91 206 -89 209
rect -75 206 -73 209
rect -65 206 -63 209
rect -55 206 -53 222
rect -29 206 -27 222
rect -19 206 -17 209
rect -2 206 0 209
rect 8 206 10 209
rect 18 206 20 209
rect 28 206 30 209
rect 44 206 46 209
rect 54 206 56 209
rect 64 206 66 222
rect 80 206 82 222
rect 90 206 92 209
rect 107 206 109 209
rect 117 206 119 209
rect 127 206 129 209
rect 137 206 139 209
rect 153 206 155 209
rect 163 206 165 209
rect 173 206 175 222
rect 189 206 191 222
rect 199 206 201 209
rect 216 206 218 209
rect 226 206 228 209
rect 236 206 238 209
rect 246 206 248 209
rect 262 206 264 209
rect 272 206 274 209
rect 282 206 284 222
rect 298 206 300 222
rect 308 206 310 209
rect 325 206 327 209
rect 335 206 337 209
rect 345 206 347 209
rect 355 206 357 209
rect 371 206 373 209
rect 381 206 383 209
rect 391 206 393 222
rect 407 206 409 222
rect 417 206 419 209
rect 434 206 436 209
rect 444 206 446 209
rect 454 206 456 209
rect 464 206 466 209
rect 480 206 482 209
rect 490 206 492 209
rect 500 206 502 222
rect 516 206 518 222
rect 526 206 528 209
rect 543 206 545 209
rect 553 206 555 209
rect 563 206 565 209
rect 573 206 575 209
rect 589 206 591 209
rect 599 206 601 209
rect 609 206 611 222
rect -257 169 -255 198
rect -247 169 -245 198
rect -230 169 -228 198
rect -220 169 -218 198
rect -210 169 -208 198
rect -200 169 -198 198
rect -184 169 -182 198
rect -174 169 -172 198
rect -164 169 -162 198
rect -148 169 -146 198
rect -138 169 -136 198
rect -121 169 -119 198
rect -111 169 -109 198
rect -101 169 -99 198
rect -91 169 -89 198
rect -75 169 -73 198
rect -65 169 -63 198
rect -55 169 -53 198
rect -29 169 -27 198
rect -19 169 -17 198
rect -2 169 0 198
rect 8 169 10 198
rect 18 169 20 198
rect 28 169 30 198
rect 44 169 46 198
rect 54 169 56 198
rect 64 169 66 198
rect 80 169 82 198
rect 90 169 92 198
rect 107 169 109 198
rect 117 169 119 198
rect 127 169 129 198
rect 137 169 139 198
rect 153 169 155 198
rect 163 169 165 198
rect 173 169 175 198
rect 189 169 191 198
rect 199 169 201 198
rect 216 169 218 198
rect 226 169 228 198
rect 236 169 238 198
rect 246 169 248 198
rect 262 169 264 198
rect 272 169 274 198
rect 282 169 284 198
rect 298 169 300 198
rect 308 169 310 198
rect 325 169 327 198
rect 335 169 337 198
rect 345 169 347 198
rect 355 169 357 198
rect 371 169 373 198
rect 381 169 383 198
rect 391 169 393 198
rect 407 169 409 198
rect 417 169 419 198
rect 434 169 436 198
rect 444 169 446 198
rect 454 169 456 198
rect 464 169 466 198
rect 480 169 482 198
rect 490 169 492 198
rect 500 169 502 198
rect 516 169 518 198
rect 526 169 528 198
rect 543 169 545 198
rect 553 169 555 198
rect 563 169 565 198
rect 573 169 575 198
rect 589 169 591 198
rect 599 169 601 198
rect 609 169 611 198
rect -257 162 -255 165
rect -247 162 -245 165
rect -230 162 -228 165
rect -220 162 -218 165
rect -210 162 -208 165
rect -200 162 -198 165
rect -184 162 -182 165
rect -174 162 -172 165
rect -164 162 -162 165
rect -148 162 -146 165
rect -138 162 -136 165
rect -121 162 -119 165
rect -111 162 -109 165
rect -332 138 -330 154
rect -322 138 -320 141
rect -305 138 -303 141
rect -295 138 -293 141
rect -285 138 -283 141
rect -275 138 -273 141
rect -259 138 -257 141
rect -249 138 -247 141
rect -239 138 -237 154
rect -223 138 -221 154
rect -213 138 -211 141
rect -196 138 -194 141
rect -186 138 -184 141
rect -176 138 -174 141
rect -166 138 -164 141
rect -150 138 -148 141
rect -140 138 -138 141
rect -130 138 -128 154
rect -114 138 -112 142
rect -101 138 -99 165
rect -91 162 -89 165
rect -75 162 -73 165
rect -65 162 -63 165
rect -55 162 -53 165
rect -29 162 -27 165
rect -19 162 -17 165
rect -2 162 0 165
rect 8 162 10 165
rect 18 155 20 165
rect 28 162 30 165
rect 44 162 46 165
rect 54 162 56 165
rect 64 162 66 165
rect 80 162 82 165
rect 90 162 92 165
rect 107 162 109 165
rect 117 162 119 165
rect 127 150 129 165
rect 137 162 139 165
rect 153 162 155 165
rect 163 162 165 165
rect 173 162 175 165
rect 189 157 191 165
rect 199 162 201 165
rect 216 162 218 165
rect 226 162 228 165
rect 236 156 238 165
rect 246 162 248 165
rect 262 162 264 165
rect 272 162 274 165
rect 282 162 284 165
rect 298 162 300 165
rect 308 162 310 165
rect 325 162 327 165
rect 335 162 337 165
rect 345 156 347 165
rect 355 162 357 165
rect 371 162 373 165
rect 381 162 383 165
rect 391 162 393 165
rect 407 162 409 165
rect 417 162 419 165
rect 434 162 436 165
rect 444 162 446 165
rect 454 156 456 165
rect 464 162 466 165
rect 480 162 482 165
rect 490 162 492 165
rect 500 162 502 165
rect 516 162 518 165
rect 526 162 528 165
rect 543 162 545 165
rect 553 162 555 165
rect 563 162 565 165
rect 573 162 575 165
rect 589 162 591 165
rect 599 162 601 165
rect 609 162 611 165
rect -83 138 -81 141
rect -73 138 -71 141
rect -54 138 -52 141
rect -34 138 -32 141
rect -10 138 -8 141
rect 0 138 2 141
rect 10 138 12 141
rect 35 138 37 142
rect 48 138 50 142
rect 66 138 68 141
rect 76 138 78 141
rect 95 138 97 141
rect 115 138 117 150
rect 139 138 141 141
rect 149 138 151 155
rect 159 138 161 141
rect 184 138 186 142
rect 197 138 199 142
rect 215 138 217 141
rect 225 138 227 141
rect 244 138 246 141
rect 264 138 266 141
rect 288 138 290 141
rect 298 138 300 141
rect 308 138 310 141
rect 333 138 335 142
rect 346 138 348 142
rect 364 138 366 141
rect 374 138 376 141
rect 390 138 392 141
rect 405 138 407 141
rect 427 138 429 141
rect 437 138 439 141
rect 447 138 449 141
rect 465 138 467 142
rect 478 138 480 142
rect 496 138 498 141
rect 506 138 508 141
rect 523 138 525 141
rect 537 138 539 141
rect 561 138 563 154
rect 571 138 573 141
rect 588 138 590 141
rect 598 138 600 141
rect 608 138 610 141
rect 618 138 620 141
rect 634 138 636 141
rect 644 138 646 141
rect 654 138 656 154
rect -332 101 -330 130
rect -322 101 -320 130
rect -305 101 -303 130
rect -295 101 -293 130
rect -285 101 -283 130
rect -275 101 -273 130
rect -259 101 -257 130
rect -249 101 -247 130
rect -239 101 -237 130
rect -223 101 -221 130
rect -213 101 -211 130
rect -196 101 -194 130
rect -186 101 -184 130
rect -176 101 -174 130
rect -166 101 -164 130
rect -150 101 -148 130
rect -140 101 -138 130
rect -130 101 -128 130
rect -332 94 -330 97
rect -322 94 -320 97
rect -305 94 -303 97
rect -295 94 -293 97
rect -285 94 -283 97
rect -275 94 -273 97
rect -259 94 -257 97
rect -249 94 -247 97
rect -239 86 -237 97
rect -223 94 -221 97
rect -213 94 -211 97
rect -196 94 -194 97
rect -186 94 -184 97
rect -176 94 -174 97
rect -166 94 -164 97
rect -150 94 -148 97
rect -140 94 -138 97
rect -130 94 -128 97
rect -114 84 -112 130
rect -101 84 -99 130
rect -83 84 -81 130
rect -73 84 -71 130
rect -54 84 -52 130
rect -34 84 -32 130
rect -114 77 -112 80
rect -101 77 -99 80
rect -83 77 -81 80
rect -73 77 -71 80
rect -54 77 -52 80
rect -34 77 -32 80
rect -10 77 -8 130
rect 0 77 2 130
rect 10 77 12 130
rect 35 84 37 130
rect 48 84 50 130
rect 66 84 68 130
rect 76 84 78 130
rect 95 84 97 130
rect 115 84 117 130
rect 35 77 37 80
rect 48 77 50 80
rect 66 77 68 80
rect 76 77 78 80
rect 95 77 97 80
rect 115 77 117 80
rect 139 77 141 130
rect 149 77 151 130
rect 159 77 161 130
rect 184 84 186 130
rect 197 84 199 130
rect 215 84 217 130
rect 225 84 227 130
rect 244 84 246 130
rect 264 84 266 130
rect 184 77 186 80
rect 197 77 199 80
rect 215 77 217 80
rect 225 77 227 80
rect 244 77 246 80
rect 264 77 266 80
rect 288 77 290 130
rect 298 77 300 130
rect 308 77 310 130
rect 333 84 335 130
rect 346 84 348 130
rect 364 84 366 130
rect 374 84 376 130
rect 390 84 392 130
rect 405 84 407 130
rect 333 77 335 80
rect 346 77 348 80
rect 364 77 366 80
rect 374 77 376 80
rect 390 77 392 80
rect 405 77 407 80
rect 427 77 429 130
rect 437 77 439 130
rect 447 77 449 130
rect 465 84 467 130
rect 478 84 480 130
rect 496 84 498 130
rect 506 84 508 130
rect 523 84 525 130
rect 537 84 539 130
rect 561 101 563 130
rect 571 101 573 130
rect 588 101 590 130
rect 598 101 600 130
rect 608 101 610 130
rect 618 101 620 130
rect 634 101 636 130
rect 644 101 646 130
rect 654 101 656 130
rect 561 94 563 97
rect 571 94 573 97
rect 588 94 590 97
rect 598 94 600 97
rect 608 88 610 97
rect 618 94 620 97
rect 634 94 636 97
rect 644 94 646 97
rect 654 94 656 97
rect 465 77 467 80
rect 478 77 480 80
rect 496 77 498 80
rect 506 77 508 80
rect 523 77 525 80
rect 537 77 539 80
rect -10 70 -8 73
rect 0 70 2 73
rect 10 70 12 73
rect 139 70 141 73
rect 149 70 151 73
rect 159 70 161 73
rect 288 70 290 73
rect 298 70 300 73
rect 308 70 310 73
rect 427 70 429 73
rect 437 70 439 73
rect 447 70 449 73
rect -279 19 -277 35
rect -269 19 -267 22
rect -252 19 -250 22
rect -242 19 -240 22
rect -232 19 -230 22
rect -222 19 -220 22
rect -206 19 -204 22
rect -196 19 -194 22
rect -186 19 -184 35
rect -170 19 -168 23
rect -157 19 -155 23
rect -139 19 -137 22
rect -129 19 -127 22
rect -110 19 -108 22
rect -90 19 -88 22
rect -66 19 -64 23
rect -53 19 -51 23
rect -35 19 -33 22
rect -25 19 -23 22
rect -6 19 -4 22
rect 14 19 16 22
rect 38 19 40 35
rect 48 19 50 35
rect 58 19 60 22
rect 88 19 90 22
rect 98 19 100 35
rect 108 19 110 22
rect 133 19 135 35
rect 143 19 145 35
rect 153 19 155 22
rect 177 19 179 35
rect 187 19 189 22
rect 197 19 199 35
rect 215 19 217 22
rect 240 19 242 22
rect 250 19 252 35
rect 260 19 262 22
rect 278 19 280 22
rect 305 19 307 22
rect 315 19 317 22
rect 325 19 327 35
rect 336 19 338 35
rect 354 19 356 22
rect 380 19 382 35
rect 390 19 392 22
rect 400 19 402 35
rect 418 19 420 22
rect 434 19 436 33
rect 444 19 446 33
rect 454 19 456 22
rect 479 19 481 22
rect 489 19 491 22
rect 499 19 501 22
rect 510 19 512 36
rect 528 19 530 22
rect 545 19 547 35
rect 555 19 557 22
rect 572 19 574 22
rect 582 19 584 22
rect 592 19 594 22
rect 602 19 604 22
rect 618 19 620 22
rect 628 19 630 22
rect 638 19 640 35
rect -279 -18 -277 11
rect -269 -18 -267 11
rect -252 -18 -250 11
rect -242 -18 -240 11
rect -232 -18 -230 11
rect -222 -18 -220 11
rect -206 -18 -204 11
rect -196 -18 -194 11
rect -186 -18 -184 11
rect -279 -25 -277 -22
rect -269 -25 -267 -22
rect -252 -25 -250 -22
rect -242 -25 -240 -22
rect -232 -31 -230 -22
rect -222 -25 -220 -22
rect -206 -25 -204 -22
rect -196 -25 -194 -22
rect -186 -25 -184 -22
rect -170 -35 -168 11
rect -157 -35 -155 11
rect -139 -35 -137 11
rect -129 -35 -127 11
rect -110 -35 -108 11
rect -90 -35 -88 11
rect -66 -35 -64 11
rect -53 -35 -51 11
rect -35 -35 -33 11
rect -25 -35 -23 11
rect -6 -35 -4 11
rect 14 -35 16 11
rect 38 -18 40 11
rect 48 -18 50 11
rect 58 -18 60 11
rect 88 -18 90 11
rect 98 -18 100 11
rect 108 -18 110 11
rect 133 -18 135 11
rect 143 -18 145 11
rect 153 -18 155 11
rect 177 -18 179 11
rect 187 -18 189 11
rect 197 -18 199 11
rect 215 -18 217 11
rect 240 -18 242 11
rect 250 -18 252 11
rect 260 -18 262 11
rect 278 -18 280 11
rect 305 -18 307 11
rect 315 -18 317 11
rect 325 -18 327 11
rect 336 -18 338 11
rect 354 -18 356 11
rect 380 -18 382 11
rect 390 -18 392 11
rect 400 -18 402 11
rect 418 -18 420 11
rect 434 -18 436 11
rect 444 -18 446 11
rect 454 -18 456 11
rect 479 -18 481 11
rect 489 -18 491 11
rect 499 -18 501 11
rect 510 -18 512 11
rect 528 -18 530 11
rect 545 -18 547 11
rect 555 -18 557 11
rect 572 -18 574 11
rect 582 -18 584 11
rect 592 -18 594 11
rect 602 -18 604 11
rect 618 -18 620 11
rect 628 -18 630 11
rect 638 -18 640 11
rect 38 -25 40 -22
rect 48 -38 50 -22
rect 58 -25 60 -22
rect 88 -25 90 -22
rect 98 -25 100 -22
rect 108 -25 110 -22
rect 133 -25 135 -22
rect 143 -25 145 -22
rect 153 -25 155 -22
rect 177 -25 179 -22
rect 187 -39 189 -22
rect 197 -39 199 -22
rect 215 -25 217 -22
rect 240 -25 242 -22
rect 250 -25 252 -22
rect 260 -25 262 -22
rect 278 -25 280 -22
rect 305 -37 307 -22
rect 315 -37 317 -22
rect 325 -25 327 -22
rect 336 -25 338 -22
rect 354 -25 356 -22
rect 380 -25 382 -22
rect 390 -37 392 -22
rect 400 -25 402 -22
rect 418 -25 420 -22
rect 434 -25 436 -22
rect 444 -25 446 -22
rect 454 -25 456 -22
rect 479 -25 481 -22
rect 489 -25 491 -22
rect 499 -33 501 -22
rect 510 -25 512 -22
rect 528 -25 530 -22
rect 545 -25 547 -22
rect 555 -25 557 -22
rect 572 -25 574 -22
rect 582 -25 584 -22
rect 592 -25 594 -22
rect 602 -25 604 -22
rect 618 -25 620 -22
rect 628 -25 630 -22
rect 638 -25 640 -22
rect -170 -42 -168 -39
rect -157 -42 -155 -39
rect -139 -42 -137 -39
rect -129 -42 -127 -39
rect -110 -42 -108 -39
rect -90 -46 -88 -39
rect -66 -42 -64 -39
rect -53 -42 -51 -39
rect -35 -42 -33 -39
rect -25 -42 -23 -39
rect -6 -42 -4 -39
rect 14 -42 16 -39
<< polycontact >>
rect -255 218 -251 222
rect -168 218 -164 222
rect -146 218 -142 222
rect -59 218 -55 222
rect -27 218 -23 222
rect 60 218 64 222
rect 82 218 86 222
rect 169 218 173 222
rect 191 218 195 222
rect 278 218 282 222
rect 300 218 304 222
rect 387 218 391 222
rect 409 218 413 222
rect 496 218 500 222
rect 518 218 522 222
rect 605 218 609 222
rect -234 185 -230 189
rect -245 178 -241 182
rect -214 185 -210 189
rect -218 172 -214 176
rect -198 185 -194 189
rect -182 171 -178 175
rect -172 184 -168 188
rect -152 185 -148 189
rect -125 185 -121 189
rect -136 178 -132 182
rect -105 185 -101 189
rect -109 172 -105 176
rect -89 185 -85 189
rect -73 171 -69 175
rect -63 184 -59 188
rect -33 185 -29 189
rect -6 185 -2 189
rect -17 178 -13 182
rect 14 185 18 189
rect 10 172 14 176
rect 30 185 34 189
rect 46 171 50 175
rect 56 184 60 188
rect 76 185 80 189
rect 103 185 107 189
rect 92 178 96 182
rect 123 185 127 189
rect 119 172 123 176
rect 139 185 143 189
rect 155 171 159 175
rect 165 184 169 188
rect 185 185 189 189
rect 212 185 216 189
rect 201 178 205 182
rect 232 185 236 189
rect 228 172 232 176
rect 248 185 252 189
rect 264 171 268 175
rect 274 184 278 188
rect 294 185 298 189
rect 321 185 325 189
rect 310 178 314 182
rect 341 185 345 189
rect 337 172 341 176
rect 357 185 361 189
rect 373 171 377 175
rect 383 184 387 188
rect 403 185 407 189
rect 430 185 434 189
rect 419 178 423 182
rect 450 185 454 189
rect 446 172 450 176
rect 466 185 470 189
rect 482 171 486 175
rect 492 184 496 188
rect 512 185 516 189
rect 539 185 543 189
rect 528 178 532 182
rect 559 185 563 189
rect 555 172 559 176
rect 575 185 579 189
rect 591 171 595 175
rect 601 184 605 188
rect -330 150 -326 154
rect -243 150 -239 154
rect -221 150 -217 154
rect -134 150 -130 154
rect 129 150 133 154
rect 145 150 149 154
rect 563 150 567 154
rect 650 150 654 154
rect -309 117 -305 121
rect -320 110 -316 114
rect -289 117 -285 121
rect -293 104 -289 108
rect -273 117 -269 121
rect -257 103 -253 107
rect -247 118 -243 122
rect -227 117 -223 121
rect -200 117 -196 121
rect -211 110 -207 114
rect -180 117 -176 121
rect -184 104 -180 108
rect -164 117 -160 121
rect -148 103 -144 107
rect -138 116 -134 120
rect -239 82 -235 86
rect -112 114 -108 118
rect -105 88 -101 92
rect -87 89 -83 93
rect -71 107 -67 111
rect -52 105 -48 109
rect -14 117 -10 121
rect -32 101 -28 105
rect -4 111 0 115
rect 6 118 10 122
rect 37 114 41 118
rect 44 88 48 92
rect 62 89 66 93
rect 78 107 82 111
rect 97 105 101 109
rect 135 117 139 121
rect 117 101 121 105
rect 145 111 149 115
rect 155 118 159 122
rect 186 114 190 118
rect 193 88 197 92
rect 211 89 215 93
rect 227 107 231 111
rect 246 105 250 109
rect 284 117 288 121
rect 266 101 270 105
rect 294 111 298 115
rect 304 118 308 122
rect 335 114 339 118
rect 342 88 346 92
rect 360 89 364 93
rect 376 107 380 111
rect 392 105 396 109
rect 423 117 427 121
rect 407 101 411 105
rect 433 111 437 115
rect 443 118 447 122
rect 467 114 471 118
rect 474 88 478 92
rect 492 89 496 93
rect 508 107 512 111
rect 525 109 529 113
rect 557 116 561 120
rect 539 109 543 113
rect 584 117 588 121
rect 573 110 577 114
rect 604 117 608 121
rect 600 104 604 108
rect 620 117 624 121
rect 636 103 640 107
rect 646 116 650 120
rect -277 31 -273 35
rect -190 31 -186 35
rect 34 31 38 35
rect 50 31 54 35
rect 100 31 104 35
rect 129 31 133 35
rect 145 31 149 35
rect 173 31 177 35
rect 199 31 203 35
rect 252 31 256 35
rect 327 31 331 35
rect 338 31 342 35
rect 376 31 380 35
rect 396 31 400 35
rect 433 33 437 37
rect 443 33 447 37
rect 506 31 510 35
rect 547 31 551 35
rect 634 31 638 35
rect -256 -2 -252 2
rect -267 -9 -263 -5
rect -236 -2 -232 2
rect -240 -15 -236 -11
rect -220 -2 -216 2
rect -204 -16 -200 -12
rect -194 -3 -190 1
rect -168 -5 -164 -1
rect -161 -31 -157 -27
rect -143 -30 -139 -26
rect -127 -12 -123 -8
rect -108 -10 -104 -6
rect -88 -10 -84 -6
rect -64 -4 -60 0
rect -57 -31 -53 -27
rect -39 -30 -35 -26
rect -23 -12 -19 -8
rect -4 -10 0 -6
rect 16 -10 20 -6
rect 54 -1 58 3
rect 84 -15 88 -11
rect 104 -9 108 -5
rect 149 -1 153 3
rect 211 -12 215 -8
rect 236 -2 240 2
rect 256 -2 260 2
rect 274 -12 278 -8
rect 350 -12 354 -8
rect 414 -12 418 -8
rect 450 -1 454 3
rect 475 -15 479 -11
rect 485 -2 489 2
rect 524 -12 528 -8
rect 541 -2 545 2
rect 568 -2 572 2
rect 557 -9 561 -5
rect 588 -2 592 2
rect 584 -15 588 -11
rect 604 -2 608 2
rect 620 -16 624 -12
rect 630 -3 634 1
rect 50 -37 54 -33
rect 183 -37 187 -33
rect 199 -37 203 -33
rect 301 -37 305 -33
rect 311 -37 315 -33
rect 386 -37 390 -33
rect 498 -37 502 -33
rect -88 -46 -84 -42
<< metal1 >>
rect -251 218 -180 221
rect -175 218 -168 221
rect -142 218 -59 221
rect -23 218 60 221
rect 86 218 169 221
rect 195 218 278 221
rect 304 218 387 221
rect 413 218 496 221
rect 522 218 605 221
rect -258 211 -243 215
rect -239 211 -216 215
rect -212 211 -170 215
rect -166 211 -153 215
rect -149 211 -134 215
rect -130 211 -107 215
rect -103 211 -61 215
rect -57 211 -34 215
rect -30 211 -15 215
rect -11 211 12 215
rect 16 211 58 215
rect 62 211 75 215
rect 79 211 94 215
rect 98 211 121 215
rect 125 211 167 215
rect 171 211 184 215
rect 188 211 203 215
rect 207 211 230 215
rect 234 211 276 215
rect 280 211 293 215
rect 297 211 312 215
rect 316 211 339 215
rect 343 211 385 215
rect 389 211 402 215
rect 406 211 421 215
rect 425 211 448 215
rect 452 211 494 215
rect 498 211 511 215
rect 515 211 530 215
rect 534 211 557 215
rect 561 211 603 215
rect 607 211 678 215
rect -262 206 -258 211
rect -240 206 -236 211
rect -216 206 -212 211
rect -193 206 -189 211
rect -170 206 -166 211
rect -153 206 -149 211
rect -131 206 -127 211
rect -107 206 -103 211
rect -84 206 -80 211
rect -61 206 -57 211
rect -34 206 -30 211
rect -12 206 -8 211
rect 12 206 16 211
rect 35 206 39 211
rect 58 206 62 211
rect 75 206 79 211
rect 97 206 101 211
rect 121 206 125 211
rect 144 206 148 211
rect 167 206 171 211
rect 184 206 188 211
rect 206 206 210 211
rect 230 206 234 211
rect 253 206 257 211
rect 276 206 280 211
rect 293 206 297 211
rect 315 206 319 211
rect 339 206 343 211
rect 362 206 366 211
rect 385 206 389 211
rect 402 206 406 211
rect 424 206 428 211
rect 448 206 452 211
rect 471 206 475 211
rect 494 206 498 211
rect 511 206 515 211
rect 533 206 537 211
rect 557 206 561 211
rect 580 206 584 211
rect 603 206 607 211
rect -253 189 -249 198
rect -226 189 -222 198
rect -206 191 -202 198
rect -253 185 -234 189
rect -226 185 -214 189
rect -253 175 -249 185
rect -241 178 -239 182
rect -226 175 -223 185
rect -205 176 -202 191
rect -180 189 -176 198
rect -194 186 -176 189
rect -161 188 -157 198
rect -144 189 -140 198
rect -117 189 -113 198
rect -97 191 -93 198
rect -194 185 -185 186
rect -262 172 -249 175
rect -262 169 -258 172
rect -235 170 -227 173
rect -214 172 -193 176
rect -235 169 -231 170
rect -197 169 -193 172
rect -189 169 -185 185
rect -168 184 -157 188
rect -154 185 -152 189
rect -144 185 -125 189
rect -117 185 -105 189
rect -179 175 -176 178
rect -178 171 -176 175
rect -161 169 -157 184
rect -144 175 -140 185
rect -132 178 -130 182
rect -153 172 -140 175
rect -117 173 -114 185
rect -96 176 -93 191
rect -71 189 -67 198
rect -85 186 -67 189
rect -52 188 -48 198
rect -25 189 -21 198
rect 2 189 6 198
rect 22 191 26 198
rect -85 185 -76 186
rect -153 169 -149 172
rect -126 170 -114 173
rect -105 172 -84 176
rect -126 169 -122 170
rect -88 169 -84 172
rect -80 169 -76 185
rect -59 184 -48 188
rect -40 185 -33 189
rect -25 185 -6 189
rect 2 185 14 189
rect -70 175 -67 178
rect -69 171 -67 175
rect -52 169 -48 184
rect -25 175 -21 185
rect -13 178 -11 182
rect 2 175 5 185
rect 23 176 26 191
rect 48 189 52 198
rect 34 186 52 189
rect 67 188 71 198
rect 84 189 88 198
rect 111 189 115 198
rect 131 191 135 198
rect 34 185 43 186
rect -34 172 -21 175
rect -34 169 -30 172
rect -7 170 1 173
rect 14 172 35 176
rect -7 169 -3 170
rect 31 169 35 172
rect 39 169 43 185
rect 60 184 71 188
rect 74 185 76 189
rect 84 185 103 189
rect 111 185 123 189
rect 49 175 52 178
rect 50 171 52 175
rect 67 169 71 184
rect 84 175 88 185
rect 96 178 98 182
rect 111 175 114 185
rect 132 176 135 191
rect 157 189 161 198
rect 143 186 161 189
rect 176 188 180 198
rect 193 189 197 198
rect 220 189 224 198
rect 240 191 244 198
rect 143 185 152 186
rect 75 172 88 175
rect 75 169 79 172
rect 102 170 110 173
rect 123 172 144 176
rect 102 169 106 170
rect 140 169 144 172
rect 148 169 152 185
rect 169 184 180 188
rect 183 185 185 189
rect 193 185 212 189
rect 220 185 232 189
rect 158 175 161 178
rect 159 171 161 175
rect 176 169 180 184
rect 193 175 197 185
rect 205 178 207 182
rect 220 175 223 185
rect 241 176 244 191
rect 266 189 270 198
rect 252 186 270 189
rect 285 188 289 198
rect 302 189 306 198
rect 329 189 333 198
rect 349 191 353 198
rect 252 185 261 186
rect 184 172 197 175
rect 184 169 188 172
rect 211 170 219 173
rect 232 172 253 176
rect 211 169 215 170
rect 249 169 253 172
rect 257 169 261 185
rect 278 184 289 188
rect 292 185 294 189
rect 302 185 321 189
rect 329 185 341 189
rect 267 175 270 178
rect 268 171 270 175
rect 285 169 289 184
rect 302 175 306 185
rect 314 178 316 182
rect 329 175 332 185
rect 350 176 353 191
rect 375 189 379 198
rect 361 186 379 189
rect 394 188 398 198
rect 411 189 415 198
rect 438 189 442 198
rect 458 191 462 198
rect 361 185 370 186
rect 293 172 306 175
rect 293 169 297 172
rect 320 170 328 173
rect 341 172 362 176
rect 320 169 324 170
rect 358 169 362 172
rect 366 169 370 185
rect 387 184 398 188
rect 401 185 403 189
rect 411 185 430 189
rect 438 185 450 189
rect 376 175 379 178
rect 377 171 379 175
rect 394 169 398 184
rect 411 175 415 185
rect 423 178 425 182
rect 438 175 441 185
rect 459 176 462 191
rect 484 189 488 198
rect 470 186 488 189
rect 503 188 507 198
rect 520 189 524 198
rect 547 189 551 198
rect 567 191 571 198
rect 470 185 479 186
rect 402 172 415 175
rect 402 169 406 172
rect 429 170 437 173
rect 450 172 471 176
rect 429 169 433 170
rect 467 169 471 172
rect 475 169 479 185
rect 496 184 507 188
rect 511 185 512 189
rect 520 185 539 189
rect 547 185 559 189
rect 485 175 488 178
rect 486 171 488 175
rect 503 169 507 184
rect 520 175 524 185
rect 532 178 534 182
rect 547 175 550 185
rect 568 176 571 191
rect 593 189 597 198
rect 579 186 597 189
rect 612 188 616 198
rect 579 185 588 186
rect 511 172 524 175
rect 511 169 515 172
rect 538 170 546 173
rect 559 172 580 176
rect 538 169 542 170
rect 576 169 580 172
rect 584 169 588 185
rect 605 184 616 188
rect 594 175 597 178
rect 595 171 597 175
rect 612 169 616 184
rect -243 161 -239 165
rect -216 161 -212 165
rect -170 161 -166 165
rect -134 161 -130 165
rect -107 161 -103 165
rect -61 161 -57 165
rect -15 161 -11 165
rect 12 161 16 165
rect 58 161 62 165
rect 94 161 98 165
rect 121 161 125 165
rect 167 161 171 165
rect 203 161 207 165
rect 230 161 234 165
rect 276 161 280 165
rect 312 161 316 165
rect 339 161 343 165
rect 385 161 389 165
rect 421 161 425 165
rect 448 161 452 165
rect 494 161 498 165
rect 530 161 534 165
rect 557 161 561 165
rect 603 161 607 165
rect -349 157 -263 161
rect -259 157 -236 161
rect -232 157 -216 161
rect -212 157 -198 161
rect -194 157 -190 161
rect -186 157 -170 161
rect -166 157 -154 161
rect -150 157 -127 161
rect -123 157 -107 161
rect -103 157 -89 161
rect -85 157 -81 161
rect -77 157 -61 161
rect -57 157 -35 161
rect -31 157 -8 161
rect -4 157 12 161
rect 16 157 30 161
rect 34 157 38 161
rect 42 157 58 161
rect 62 157 74 161
rect 78 157 101 161
rect 105 157 121 161
rect 125 157 139 161
rect 143 157 147 161
rect 151 157 167 161
rect 171 157 183 161
rect 187 157 210 161
rect 214 157 230 161
rect 234 157 248 161
rect 252 157 256 161
rect 260 157 276 161
rect 280 157 292 161
rect 296 157 319 161
rect 323 157 339 161
rect 343 157 357 161
rect 361 157 365 161
rect 369 157 385 161
rect 389 157 401 161
rect 405 157 428 161
rect 432 157 448 161
rect 452 157 466 161
rect 470 157 474 161
rect 478 157 494 161
rect 498 157 510 161
rect 514 157 537 161
rect 541 157 557 161
rect 561 157 575 161
rect 579 157 583 161
rect 587 157 603 161
rect -349 93 -345 157
rect -326 150 -243 153
rect -217 150 -134 153
rect 133 150 145 154
rect 567 150 650 153
rect 674 147 678 211
rect -333 143 -318 147
rect -314 143 -291 147
rect -287 143 -245 147
rect -241 143 -228 147
rect -224 143 -209 147
rect -205 143 -182 147
rect -178 143 -136 147
rect -132 143 -121 147
rect -117 143 -96 147
rect -92 143 -88 147
rect -84 143 -69 147
rect -65 143 -28 147
rect -24 143 -15 147
rect -11 143 14 147
rect 18 143 28 147
rect 32 143 53 147
rect 57 143 61 147
rect 65 143 80 147
rect 84 143 121 147
rect 125 143 134 147
rect 138 143 163 147
rect 167 143 177 147
rect 181 143 202 147
rect 206 143 210 147
rect 214 143 229 147
rect 233 143 270 147
rect 274 143 283 147
rect 287 143 312 147
rect 316 143 326 147
rect 330 143 351 147
rect 355 143 359 147
rect 363 143 378 147
rect 382 143 411 147
rect 415 143 422 147
rect 426 143 451 147
rect 455 143 467 147
rect 471 143 483 147
rect 487 143 491 147
rect 495 143 510 147
rect 514 143 543 147
rect 547 143 556 147
rect 560 143 575 147
rect 579 143 602 147
rect 606 143 648 147
rect 652 143 678 147
rect -337 138 -333 143
rect -315 138 -311 143
rect -291 138 -287 143
rect -268 138 -264 143
rect -245 138 -241 143
rect -228 138 -224 143
rect -206 138 -202 143
rect -182 138 -178 143
rect -159 138 -155 143
rect -136 138 -132 143
rect -106 138 -102 143
rect -69 138 -65 143
rect -15 138 -11 143
rect 4 138 8 143
rect 43 138 47 143
rect 80 138 84 143
rect 134 138 138 143
rect 153 138 157 143
rect 192 138 196 143
rect 229 138 233 143
rect 283 138 287 143
rect 302 138 306 143
rect 341 138 345 143
rect 378 138 382 143
rect 422 138 426 143
rect 441 138 445 143
rect 473 138 477 143
rect 510 138 514 143
rect 556 138 560 143
rect 578 138 582 143
rect 602 138 606 143
rect 625 138 629 143
rect 648 138 652 143
rect -328 121 -324 130
rect -301 121 -297 130
rect -281 123 -277 130
rect -328 117 -309 121
rect -301 117 -289 121
rect -328 107 -324 117
rect -316 110 -314 114
rect -301 107 -298 117
rect -280 108 -277 123
rect -255 121 -251 130
rect -236 122 -232 130
rect -269 118 -251 121
rect -243 118 -232 122
rect -219 121 -215 130
rect -192 123 -188 130
rect -172 123 -168 130
rect -269 117 -260 118
rect -337 104 -324 107
rect -337 101 -333 104
rect -310 102 -302 105
rect -289 104 -268 108
rect -310 101 -306 102
rect -272 101 -268 104
rect -264 101 -260 117
rect -254 107 -251 110
rect -253 103 -251 107
rect -236 101 -232 118
rect -229 117 -227 121
rect -219 117 -200 121
rect -188 118 -180 121
rect -192 117 -180 118
rect -219 107 -215 117
rect -207 110 -205 114
rect -228 104 -215 107
rect -192 105 -189 117
rect -171 108 -168 123
rect -146 121 -142 130
rect -160 118 -142 121
rect -127 120 -123 130
rect -160 117 -151 118
rect -228 101 -224 104
rect -201 102 -189 105
rect -180 104 -159 108
rect -201 101 -197 102
rect -163 101 -159 104
rect -155 101 -151 117
rect -134 116 -123 120
rect -145 107 -142 110
rect -144 103 -142 107
rect -127 101 -123 116
rect -318 93 -314 97
rect -291 93 -287 97
rect -245 93 -241 97
rect -209 93 -205 97
rect -182 93 -178 97
rect -136 93 -132 97
rect -349 89 -338 93
rect -334 89 -311 93
rect -307 89 -291 93
rect -287 89 -273 93
rect -269 89 -265 93
rect -261 89 -245 93
rect -241 89 -229 93
rect -225 89 -202 93
rect -198 89 -182 93
rect -178 89 -164 93
rect -160 89 -156 93
rect -152 89 -136 93
rect -301 -26 -297 89
rect -239 75 -236 82
rect -136 69 -132 89
rect -119 90 -115 130
rect -108 114 -107 118
rect -98 93 -94 130
rect -88 121 -84 130
rect -31 121 -27 130
rect -6 122 -2 130
rect -88 116 -27 121
rect -79 112 -75 116
rect -18 117 -14 120
rect -6 118 6 122
rect -67 107 -66 111
rect -122 86 -115 90
rect -106 88 -105 92
rect -98 89 -87 93
rect -119 84 -115 86
rect -98 84 -94 89
rect -79 84 -75 107
rect -48 105 -44 109
rect -7 105 -4 115
rect -28 101 -24 105
rect -19 101 -4 105
rect -69 87 -27 91
rect -69 84 -65 87
rect -31 84 -27 87
rect 4 84 8 118
rect -109 69 -105 80
rect -88 76 -84 80
rect -69 76 -65 80
rect -88 72 -65 76
rect -15 80 8 84
rect 13 84 17 130
rect 30 90 34 130
rect 41 114 42 118
rect 51 93 55 130
rect 61 121 65 130
rect 118 121 122 130
rect 143 122 147 130
rect 61 116 122 121
rect 70 112 74 116
rect 131 117 135 120
rect 143 118 155 122
rect 82 107 83 111
rect 27 86 34 90
rect 43 88 44 92
rect 51 89 62 93
rect 30 84 34 86
rect 51 84 55 89
rect 70 84 74 107
rect 101 105 105 109
rect 142 105 145 115
rect 121 101 125 105
rect 130 101 145 105
rect -50 69 -46 80
rect -15 77 -11 80
rect 80 87 122 91
rect 80 84 84 87
rect 118 84 122 87
rect 153 84 157 118
rect 13 77 17 79
rect 4 69 8 73
rect 40 69 44 80
rect 61 76 65 80
rect 80 76 84 80
rect 61 72 84 76
rect 134 80 157 84
rect 162 86 166 130
rect 179 95 183 130
rect 190 114 191 118
rect 176 91 183 95
rect 200 93 204 130
rect 210 121 214 130
rect 267 121 271 130
rect 292 122 296 130
rect 210 116 271 121
rect 219 112 223 116
rect 280 117 284 120
rect 292 118 304 122
rect 231 107 232 111
rect 179 84 183 91
rect 192 88 193 92
rect 200 89 211 93
rect 200 84 204 89
rect 219 84 223 107
rect 250 105 254 109
rect 291 105 294 115
rect 270 101 274 105
rect 279 101 294 105
rect 99 69 103 80
rect 134 77 138 80
rect 162 77 166 81
rect 229 87 271 91
rect 229 84 233 87
rect 267 84 271 87
rect 302 84 306 118
rect 153 69 157 73
rect 189 69 193 80
rect 210 76 214 80
rect 229 76 233 80
rect 210 72 233 76
rect 283 80 306 84
rect 311 113 315 130
rect 311 110 317 113
rect 311 85 315 110
rect 328 95 332 130
rect 339 114 340 118
rect 325 91 332 95
rect 349 93 353 130
rect 359 121 363 130
rect 408 121 412 130
rect 431 122 435 130
rect 359 116 412 121
rect 368 112 372 116
rect 421 117 423 120
rect 431 118 443 122
rect 380 107 381 111
rect 328 84 332 91
rect 341 88 342 92
rect 349 89 360 93
rect 349 84 353 89
rect 368 84 372 107
rect 396 105 399 109
rect 430 105 433 115
rect 411 101 415 105
rect 420 101 433 105
rect 378 87 412 91
rect 378 84 382 87
rect 408 84 412 87
rect 441 84 445 118
rect 248 69 252 80
rect 283 77 287 80
rect 311 77 315 80
rect 302 69 306 73
rect 338 69 342 80
rect 359 76 363 80
rect 378 76 382 80
rect 359 72 382 76
rect 422 80 445 84
rect 450 82 454 130
rect 460 104 464 130
rect 471 114 472 118
rect 460 84 464 99
rect 481 93 485 130
rect 491 121 495 130
rect 540 121 544 130
rect 491 120 544 121
rect 565 121 569 130
rect 592 121 596 130
rect 612 123 616 130
rect 491 116 557 120
rect 565 117 584 121
rect 592 117 604 121
rect 500 112 504 116
rect 512 107 513 111
rect 529 109 531 113
rect 543 109 544 113
rect 565 107 569 117
rect 577 110 579 114
rect 592 107 595 117
rect 613 108 616 123
rect 638 121 642 130
rect 624 118 642 121
rect 657 120 661 130
rect 624 117 633 118
rect 473 88 474 92
rect 481 89 492 93
rect 481 84 485 89
rect 500 84 504 107
rect 556 104 569 107
rect 556 101 560 104
rect 583 102 591 105
rect 604 104 625 108
rect 583 101 587 102
rect 621 101 625 104
rect 629 101 633 117
rect 650 116 661 120
rect 639 107 642 110
rect 640 103 642 107
rect 657 101 661 116
rect 575 93 579 97
rect 602 93 606 97
rect 648 93 652 97
rect 394 69 398 80
rect 422 77 426 80
rect 510 87 544 91
rect 510 84 514 87
rect 540 84 544 87
rect 441 69 445 73
rect 470 69 474 80
rect 491 76 495 80
rect 510 76 514 80
rect 491 72 514 76
rect 559 89 582 93
rect 586 89 602 93
rect 606 89 620 93
rect 624 89 628 93
rect 632 89 648 93
rect 527 69 531 80
rect 555 69 559 89
rect -136 65 -125 69
rect -121 65 -107 69
rect -103 65 -89 69
rect -85 65 -56 69
rect -52 65 -26 69
rect -22 65 -16 69
rect -12 65 13 69
rect 17 65 24 69
rect 28 65 42 69
rect 46 65 60 69
rect 64 65 93 69
rect 97 65 123 69
rect 127 65 133 69
rect 137 65 162 69
rect 166 65 173 69
rect 177 65 191 69
rect 195 65 209 69
rect 213 65 242 69
rect 246 65 272 69
rect 276 65 282 69
rect 286 65 311 69
rect 315 65 322 69
rect 326 65 340 69
rect 344 65 358 69
rect 362 65 388 69
rect 392 65 413 69
rect 417 65 421 69
rect 425 65 450 69
rect 454 65 458 69
rect 462 65 472 69
rect 476 65 490 69
rect 494 65 523 69
rect 527 65 555 69
rect -273 31 -200 34
rect 13 35 18 41
rect 57 35 60 56
rect 186 54 189 57
rect 111 35 116 49
rect 146 51 203 54
rect 146 35 149 51
rect 174 35 177 41
rect 200 35 203 51
rect 312 38 315 57
rect 358 46 361 57
rect 358 41 360 46
rect -195 31 -190 34
rect 13 31 34 35
rect 54 31 60 35
rect 104 31 129 35
rect 256 33 312 34
rect 328 35 331 41
rect 256 31 317 33
rect 358 34 361 41
rect 396 35 399 50
rect 424 43 447 46
rect 342 31 376 34
rect 444 37 447 43
rect 424 34 433 37
rect 437 34 439 37
rect 503 31 506 34
rect 551 31 634 34
rect 674 28 678 143
rect -280 24 -265 28
rect -261 24 -238 28
rect -234 24 -192 28
rect -188 24 -177 28
rect -173 24 -152 28
rect -148 24 -144 28
rect -140 24 -125 28
rect -121 24 -84 28
rect -80 24 -73 28
rect -69 24 -48 28
rect -44 24 -40 28
rect -36 24 -21 28
rect -17 24 20 28
rect 24 24 33 28
rect 37 24 62 28
rect 66 24 83 28
rect 87 24 112 28
rect 116 24 128 28
rect 132 24 157 28
rect 161 24 172 28
rect 176 24 201 28
rect 205 24 220 28
rect 224 24 235 28
rect 239 24 264 28
rect 268 24 283 28
rect 287 24 300 28
rect 304 24 331 28
rect 335 24 359 28
rect 363 24 375 28
rect 379 24 404 28
rect 408 24 429 28
rect 433 24 458 28
rect 462 24 474 28
rect 478 24 505 28
rect 509 24 540 28
rect 544 24 559 28
rect 563 24 586 28
rect 590 24 632 28
rect 636 24 678 28
rect -284 19 -280 24
rect -262 19 -258 24
rect -238 19 -234 24
rect -215 19 -211 24
rect -192 19 -188 24
rect -162 19 -158 24
rect -125 19 -121 24
rect -58 19 -54 24
rect -21 19 -17 24
rect 33 19 37 24
rect 52 19 56 24
rect 102 19 106 24
rect 128 19 132 24
rect 147 19 151 24
rect 172 19 176 24
rect 191 19 195 24
rect 210 19 214 24
rect 235 19 239 24
rect 273 19 277 24
rect 300 19 304 24
rect 319 19 323 24
rect 339 19 343 24
rect -275 2 -271 11
rect -248 2 -244 11
rect -228 4 -224 11
rect -275 -2 -256 2
rect -248 -2 -236 2
rect -275 -12 -271 -2
rect -263 -9 -261 -5
rect -248 -12 -245 -2
rect -227 -11 -224 4
rect -202 2 -198 11
rect -216 -1 -198 2
rect -183 1 -179 11
rect -216 -2 -207 -1
rect -284 -15 -271 -12
rect -284 -18 -280 -15
rect -257 -17 -249 -14
rect -236 -15 -215 -11
rect -257 -18 -253 -17
rect -219 -18 -215 -15
rect -211 -18 -207 -2
rect -190 -3 -179 1
rect -201 -12 -198 -9
rect -200 -16 -198 -12
rect -183 -18 -179 -3
rect -175 -15 -171 11
rect -164 -5 -163 -1
rect -265 -26 -261 -22
rect -238 -26 -234 -22
rect -192 -26 -188 -22
rect -301 -30 -285 -26
rect -281 -30 -258 -26
rect -254 -30 -238 -26
rect -234 -30 -220 -26
rect -216 -30 -212 -26
rect -208 -30 -192 -26
rect -192 -50 -188 -30
rect -175 -35 -171 -20
rect -154 -26 -150 11
rect -144 2 -140 11
rect -87 2 -83 11
rect -144 -3 -83 2
rect -135 -7 -131 -3
rect -123 -12 -122 -8
rect -104 -10 -100 -6
rect -84 -10 -80 -6
rect -162 -31 -161 -27
rect -154 -30 -143 -26
rect -154 -35 -150 -30
rect -135 -35 -131 -12
rect -71 -15 -67 11
rect -60 -4 -59 0
rect -125 -32 -83 -28
rect -125 -35 -121 -32
rect -87 -35 -83 -32
rect -165 -50 -161 -39
rect -144 -43 -140 -39
rect -125 -43 -121 -39
rect -144 -47 -121 -43
rect -71 -35 -67 -20
rect -50 -26 -46 11
rect -40 2 -36 11
rect 17 2 21 11
rect -40 -3 21 2
rect 42 3 46 11
rect 42 -1 54 3
rect -31 -7 -27 -3
rect -19 -12 -18 -8
rect 0 -10 4 -7
rect 20 -10 24 -6
rect 52 -11 56 -1
rect -58 -31 -57 -27
rect -50 -30 -39 -26
rect -50 -35 -46 -30
rect -31 -35 -27 -12
rect 33 -15 56 -11
rect 61 -12 65 11
rect 349 19 353 24
rect 375 19 379 24
rect 394 19 398 24
rect 413 19 417 24
rect 429 19 433 24
rect 448 19 452 24
rect 474 19 478 24
rect 523 19 527 24
rect 540 19 544 24
rect 562 19 566 24
rect 586 19 590 24
rect 609 19 613 24
rect 632 19 636 24
rect 83 -5 87 11
rect 83 -8 104 -5
rect 61 -15 84 -12
rect 33 -18 37 -15
rect 61 -18 65 -15
rect 92 -18 96 -8
rect 111 -6 115 11
rect 137 3 141 11
rect 137 -1 149 3
rect 147 -11 151 -1
rect 111 -18 115 -11
rect 128 -15 151 -11
rect 156 -10 160 11
rect 181 3 185 11
rect 200 3 204 11
rect 181 -1 204 3
rect 200 -8 204 -1
rect 218 -6 222 11
rect 230 -2 236 1
rect 254 -2 256 2
rect 254 -6 257 -2
rect 156 -15 159 -10
rect 200 -12 211 -8
rect 218 -9 257 -6
rect 263 -8 267 11
rect 128 -18 132 -15
rect 156 -18 160 -15
rect 200 -18 204 -12
rect 218 -18 222 -9
rect 263 -12 274 -8
rect 244 -15 267 -12
rect 244 -18 248 -15
rect 263 -18 267 -15
rect 281 -18 285 11
rect 309 -1 313 11
rect 329 -1 333 11
rect 309 -4 343 -1
rect 339 -8 343 -4
rect 339 -12 350 -8
rect 339 -18 343 -12
rect 357 -18 361 11
rect 384 3 388 11
rect 403 3 407 11
rect 384 -1 407 3
rect 403 -8 407 -1
rect 403 -12 414 -8
rect 421 -9 425 11
rect 438 3 442 11
rect 438 -1 450 3
rect 403 -18 407 -12
rect 448 -11 452 -1
rect 421 -18 425 -14
rect 429 -15 452 -11
rect 457 -11 461 11
rect 476 -2 485 1
rect 513 -8 517 11
rect 531 2 535 11
rect 549 2 553 11
rect 576 2 580 11
rect 596 4 600 11
rect 531 -2 541 2
rect 549 -2 568 2
rect 576 -2 588 2
rect 457 -15 475 -11
rect 513 -12 524 -8
rect 483 -15 517 -12
rect 429 -18 433 -15
rect 457 -18 461 -15
rect 483 -18 487 -15
rect 504 -18 508 -15
rect 531 -18 535 -2
rect 549 -12 553 -2
rect 561 -9 563 -5
rect 576 -12 579 -2
rect 597 -11 600 4
rect 622 2 626 11
rect 608 -1 626 2
rect 641 1 645 11
rect 608 -2 617 -1
rect 52 -26 56 -22
rect 83 -26 87 -22
rect 102 -26 106 -22
rect 147 -26 151 -22
rect 172 -26 176 -22
rect 210 -26 214 -22
rect 235 -26 239 -22
rect 254 -26 258 -22
rect 273 -26 277 -22
rect 300 -26 304 -22
rect 349 -26 353 -22
rect 375 -26 379 -22
rect 413 -26 417 -22
rect 448 -26 452 -22
rect 474 -26 478 -22
rect 493 -26 497 -22
rect 513 -26 517 -22
rect 540 -15 553 -12
rect 540 -18 544 -15
rect 567 -17 575 -14
rect 588 -15 609 -11
rect 567 -18 571 -17
rect 605 -18 609 -15
rect 613 -18 617 -2
rect 634 -3 645 1
rect 623 -12 626 -9
rect 624 -16 626 -12
rect 641 -18 645 -3
rect 523 -26 527 -22
rect 559 -26 563 -22
rect 586 -26 590 -22
rect 632 -26 636 -22
rect -21 -32 21 -28
rect -21 -35 -17 -32
rect 17 -35 21 -32
rect -106 -50 -102 -39
rect -84 -46 -82 -42
rect -61 -50 -57 -39
rect -40 -43 -36 -39
rect -21 -43 -17 -39
rect -40 -47 -17 -43
rect 36 -30 61 -26
rect 65 -30 82 -26
rect 86 -30 111 -26
rect 115 -30 127 -26
rect 131 -30 156 -26
rect 160 -30 171 -26
rect 175 -30 200 -26
rect 204 -30 222 -26
rect 226 -30 235 -26
rect 239 -30 263 -26
rect 267 -30 285 -26
rect 289 -30 300 -26
rect 304 -30 330 -26
rect 334 -30 361 -26
rect 365 -30 374 -26
rect 378 -30 403 -26
rect 407 -30 425 -26
rect 429 -30 433 -26
rect 437 -30 457 -26
rect 461 -30 474 -26
rect 478 -30 504 -26
rect 508 -30 535 -26
rect 543 -30 566 -26
rect 570 -30 586 -26
rect 590 -30 604 -26
rect 608 -30 612 -26
rect 616 -30 632 -26
rect -2 -50 2 -39
rect 32 -50 36 -30
rect 54 -37 183 -34
rect 203 -34 301 -33
rect 203 -36 293 -34
rect 59 -42 64 -37
rect 184 -42 187 -37
rect 298 -36 301 -34
rect 312 -42 315 -37
rect 383 -37 386 -34
rect 495 -37 498 -34
rect 184 -45 315 -42
rect -188 -54 -163 -50
rect -159 -54 -145 -50
rect -141 -54 -112 -50
rect -108 -54 -82 -50
rect -78 -54 -61 -50
rect -57 -54 -41 -50
rect -37 -54 -8 -50
rect -4 -54 22 -50
rect 26 -54 36 -50
<< m2contact >>
rect -180 218 -175 223
rect -239 177 -234 182
rect -227 170 -222 175
rect -180 178 -175 183
rect -130 177 -125 182
rect -71 178 -66 183
rect -11 177 -6 182
rect 1 170 6 175
rect 48 178 53 183
rect 98 177 103 182
rect 110 170 115 175
rect 157 178 162 183
rect 207 177 212 182
rect 219 170 224 175
rect 266 178 271 183
rect 316 177 321 182
rect 328 170 333 175
rect 375 178 380 183
rect 425 177 430 182
rect 437 170 442 175
rect 484 178 489 183
rect 534 177 539 182
rect 546 170 551 175
rect 593 178 598 183
rect -314 109 -309 114
rect -302 102 -297 107
rect -254 110 -249 115
rect -193 118 -188 123
rect -205 109 -200 114
rect -146 110 -141 115
rect -239 70 -234 75
rect -127 86 -122 91
rect -107 114 -102 119
rect -23 115 -18 120
rect -79 107 -74 112
rect -66 107 -61 112
rect -111 88 -106 93
rect -44 104 -39 109
rect -24 100 -19 105
rect 22 86 27 91
rect 42 114 47 119
rect 126 115 131 120
rect 70 107 75 112
rect 83 107 88 112
rect 38 88 43 93
rect 105 104 110 109
rect 125 100 130 105
rect 13 79 18 84
rect 171 91 176 96
rect 191 114 196 119
rect 275 115 280 120
rect 219 107 224 112
rect 232 107 237 112
rect 162 81 167 86
rect 187 88 192 93
rect 254 104 259 109
rect 274 100 279 105
rect 320 91 325 96
rect 340 114 345 119
rect 416 115 421 120
rect 368 107 373 112
rect 381 107 386 112
rect 311 80 316 85
rect 336 88 341 93
rect 399 104 404 109
rect 415 100 420 105
rect 472 114 477 119
rect 460 99 465 104
rect 500 107 505 112
rect 513 107 518 112
rect 531 108 536 113
rect 544 108 549 113
rect 579 109 584 114
rect 591 102 596 107
rect 638 110 643 115
rect 450 77 455 82
rect 56 56 61 61
rect 186 57 191 62
rect 311 57 316 62
rect 357 57 362 62
rect -200 31 -195 36
rect 111 49 116 54
rect 174 41 179 46
rect 396 50 401 55
rect 327 41 332 46
rect 360 41 365 46
rect 312 33 317 38
rect 419 42 424 47
rect 419 33 424 38
rect 498 31 503 36
rect -261 -10 -256 -5
rect -249 -17 -244 -12
rect -202 -9 -197 -4
rect -163 -5 -158 0
rect -175 -20 -170 -15
rect -135 -12 -130 -7
rect -122 -12 -117 -7
rect -100 -11 -95 -6
rect -80 -11 -75 -6
rect -167 -31 -162 -26
rect -59 -4 -54 1
rect -72 -20 -67 -15
rect -31 -12 -26 -7
rect -18 -12 -13 -7
rect 4 -11 9 -6
rect 24 -11 29 -6
rect -63 -31 -58 -26
rect 111 -11 116 -6
rect 225 -2 230 3
rect 159 -15 164 -10
rect 361 -3 366 2
rect 421 -14 426 -9
rect 471 -3 476 2
rect 563 -10 568 -5
rect 575 -17 580 -12
rect 622 -9 627 -4
rect -82 -47 -77 -42
rect 59 -47 64 -42
rect 293 -39 298 -34
rect 378 -38 383 -33
rect 490 -39 495 -34
<< metal2 >>
rect -180 203 -177 218
rect -180 200 -137 203
rect -262 179 -239 182
rect -254 115 -251 179
rect -234 179 -180 182
rect -175 179 -130 182
rect -125 179 -71 182
rect -66 179 -11 182
rect -6 179 48 182
rect 53 179 98 182
rect 103 179 157 182
rect 162 179 207 182
rect 212 179 266 182
rect 271 179 316 182
rect 321 179 375 182
rect 380 179 425 182
rect 430 179 484 182
rect 489 179 534 182
rect 539 179 593 182
rect -222 171 -166 174
rect -188 119 -115 122
rect -119 116 -107 119
rect -309 111 -254 114
rect -312 102 -302 105
rect -261 -5 -258 111
rect -249 111 -205 114
rect -200 111 -146 114
rect -102 116 -23 119
rect -63 115 -23 116
rect 2 119 5 170
rect 2 116 42 119
rect -63 112 -59 115
rect 47 116 126 119
rect 86 115 126 116
rect 220 119 223 170
rect 329 155 332 170
rect 289 152 332 155
rect 438 153 441 170
rect 547 153 550 170
rect 86 112 90 115
rect 196 116 275 119
rect 235 115 275 116
rect 235 112 239 115
rect -130 107 -79 110
rect -61 107 -59 112
rect 62 107 70 110
rect 88 107 90 112
rect -44 103 -40 104
rect -126 100 -40 103
rect 211 107 219 110
rect 237 107 239 112
rect 105 100 109 104
rect -126 91 -123 100
rect -24 91 -21 100
rect 23 97 109 100
rect 254 103 258 104
rect 172 100 258 103
rect 289 104 292 152
rect 353 150 441 153
rect 478 150 550 153
rect 353 135 356 150
rect 478 136 481 150
rect 341 132 356 135
rect 440 133 481 136
rect 341 119 344 132
rect 345 116 416 119
rect 384 115 416 116
rect 384 112 388 115
rect 361 108 368 111
rect 386 107 388 112
rect 279 101 292 104
rect 398 104 399 107
rect 398 103 402 104
rect 321 100 402 103
rect 440 104 443 133
rect 460 116 472 119
rect 477 116 520 119
rect 516 112 520 116
rect 594 114 597 178
rect 491 107 500 110
rect 518 107 520 112
rect 584 111 638 114
rect 420 101 443 104
rect 23 91 26 97
rect -106 88 -21 91
rect -102 76 -99 88
rect 125 91 128 100
rect 172 96 175 100
rect 43 88 128 91
rect 275 91 278 100
rect 321 96 324 100
rect 192 88 278 91
rect 415 91 418 100
rect 531 103 534 108
rect 465 100 534 103
rect 341 88 418 91
rect 545 91 548 108
rect 473 88 548 91
rect -234 70 -173 73
rect -117 73 -99 76
rect -206 31 -200 34
rect -163 0 -159 41
rect -58 1 -55 57
rect 13 46 18 79
rect 47 76 50 88
rect 34 73 50 76
rect 57 61 60 71
rect 163 53 166 81
rect 196 76 199 88
rect 180 73 199 76
rect 312 62 315 80
rect 345 76 348 88
rect 357 76 360 77
rect 331 73 348 76
rect 357 62 360 71
rect 191 58 195 61
rect 116 50 396 53
rect 18 42 174 45
rect 179 42 327 45
rect 365 43 419 46
rect 317 34 419 37
rect 451 34 454 77
rect 451 31 498 34
rect -256 -8 -202 -5
rect -158 -3 -115 0
rect -119 -7 -115 -3
rect -54 -3 -11 0
rect -143 -12 -135 -9
rect -117 -12 -115 -7
rect -15 -7 -11 -3
rect 160 -2 225 1
rect -244 -16 -213 -13
rect -100 -16 -97 -11
rect -170 -19 -97 -16
rect -80 -28 -77 -11
rect -38 -12 -31 -9
rect -13 -12 -11 -7
rect 29 -10 111 -7
rect 160 -10 163 -2
rect 366 -3 471 0
rect 580 -5 583 109
rect 596 103 667 106
rect 5 -16 8 -11
rect -67 -19 8 -16
rect -162 -31 -77 -28
rect 24 -28 27 -11
rect 568 -8 622 -5
rect -58 -31 27 -28
rect 298 -37 378 -34
rect 422 -34 425 -14
rect 580 -16 651 -13
rect 422 -37 490 -34
rect -77 -46 59 -43
<< m3contact >>
rect -137 199 -132 204
rect -135 106 -130 111
rect 57 106 62 111
rect 206 107 211 112
rect 356 107 361 112
rect 455 115 460 120
rect -173 69 -168 74
rect -59 57 -54 62
rect -164 41 -158 46
rect -211 30 -206 35
rect 56 71 61 76
rect 356 71 361 76
rect 195 57 200 62
rect -148 -12 -143 -7
rect -43 -12 -38 -7
<< m123contact >>
rect 468 88 473 93
rect 13 41 18 46
rect 285 -7 290 -2
<< metal3 >>
rect -138 204 -131 205
rect -138 199 -137 204
rect -132 199 -131 204
rect -138 198 -131 199
rect -136 112 -133 198
rect 205 112 212 113
rect -136 111 -129 112
rect -136 106 -135 111
rect -130 106 -129 111
rect -136 105 -129 106
rect 56 111 63 112
rect 56 106 57 111
rect 62 106 63 111
rect 205 107 206 112
rect 211 107 212 112
rect 456 111 459 115
rect 361 108 459 111
rect 205 106 212 107
rect 56 105 63 106
rect 57 76 60 105
rect -174 74 -167 75
rect -174 69 -173 74
rect -168 69 -167 74
rect -174 68 -167 69
rect -172 62 -169 68
rect 194 62 201 63
rect 194 61 195 62
rect -54 58 195 61
rect 194 57 195 58
rect 200 61 201 62
rect 209 61 212 106
rect 357 76 360 107
rect 200 58 212 61
rect 200 57 201 58
rect 194 56 201 57
rect -158 42 13 45
rect -212 35 -205 36
rect -212 30 -211 35
rect -206 34 -205 35
rect -206 31 -144 34
rect -206 30 -205 31
rect -212 29 -205 30
rect -147 -6 -144 31
rect -42 -6 -39 32
rect -149 -7 -142 -6
rect -149 -12 -148 -7
rect -143 -12 -142 -7
rect -149 -13 -142 -12
rect -44 -7 -37 -6
rect 469 -3 472 88
rect 290 -6 472 -3
rect -44 -12 -43 -7
rect -38 -12 -37 -7
rect -44 -13 -37 -12
<< m4contact >>
rect -172 57 -167 62
rect -42 32 -37 37
<< metal4 >>
rect -172 53 -169 57
rect -172 50 -38 53
rect -41 37 -38 50
<< labels >>
rlabel metal1 99 145 99 145 5 vdd
rlabel metal1 79 67 79 67 1 gnd
rlabel metal1 317 110 317 113 1 g2
rlabel metal1 15 93 15 98 1 c1
rlabel m2contact 358 58 361 58 1 p3
rlabel m2contact 113 54 116 54 6 g1
rlabel metal1 282 -5 284 -5 1 c3
rlabel metal1 113 -3 115 -3 1 c2
rlabel space 311 55 315 55 6 g2
rlabel metal1 -40 185 -40 189 1 b1
rlabel metal1 511 185 511 189 1 a3
rlabel metal1 401 185 401 189 1 b3
rlabel metal1 292 185 292 189 1 a2
rlabel metal1 183 185 183 189 1 b2
rlabel metal1 74 185 74 189 1 a1
rlabel metal2 667 103 667 106 7 sum3
rlabel metal2 -262 179 -262 182 3 clk
rlabel metal2 -166 171 -166 174 1 sum0
rlabel metal1 -154 185 -154 189 1 a0
rlabel metal2 651 -16 651 -13 1 c4
rlabel metal2 -213 -16 -213 -13 1 sum1
rlabel metal1 -229 117 -229 121 1 b0
rlabel metal2 -312 102 -312 105 1 sum2
<< end >>
