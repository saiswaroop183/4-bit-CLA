magic
tech scmos
timestamp 1638628949
<< nwell >>
rect 32 -3 558 24
<< ntransistor >>
rect 43 -29 45 -25
rect 53 -29 55 -25
rect 63 -29 65 -25
rect 93 -29 95 -25
rect 103 -29 105 -25
rect 113 -29 115 -25
rect 138 -29 140 -25
rect 148 -29 150 -25
rect 158 -29 160 -25
rect 182 -29 184 -25
rect 192 -29 194 -25
rect 202 -29 204 -25
rect 220 -29 222 -25
rect 245 -29 247 -25
rect 255 -29 257 -25
rect 265 -29 267 -25
rect 283 -29 285 -25
rect 310 -29 312 -25
rect 320 -29 322 -25
rect 330 -29 332 -25
rect 341 -29 343 -25
rect 359 -29 361 -25
rect 385 -29 387 -25
rect 395 -29 397 -25
rect 405 -29 407 -25
rect 423 -29 425 -25
rect 449 -29 451 -25
rect 459 -29 461 -25
rect 469 -29 471 -25
rect 494 -29 496 -25
rect 504 -29 506 -25
rect 514 -29 516 -25
rect 525 -29 527 -25
rect 543 -29 545 -25
<< ptransistor >>
rect 43 4 45 12
rect 53 4 55 12
rect 63 4 65 12
rect 93 4 95 12
rect 103 4 105 12
rect 113 4 115 12
rect 138 4 140 12
rect 148 4 150 12
rect 158 4 160 12
rect 182 4 184 12
rect 192 4 194 12
rect 202 4 204 12
rect 220 4 222 12
rect 245 4 247 12
rect 255 4 257 12
rect 265 4 267 12
rect 283 4 285 12
rect 310 4 312 12
rect 320 4 322 12
rect 330 4 332 12
rect 341 4 343 12
rect 359 4 361 12
rect 385 4 387 12
rect 395 4 397 12
rect 405 4 407 12
rect 423 4 425 12
rect 449 4 451 12
rect 459 4 461 12
rect 469 4 471 12
rect 494 4 496 12
rect 504 4 506 12
rect 514 4 516 12
rect 525 4 527 12
rect 543 4 545 12
<< ndiffusion >>
rect 42 -29 43 -25
rect 45 -29 53 -25
rect 55 -29 57 -25
rect 61 -29 63 -25
rect 65 -29 66 -25
rect 92 -29 93 -25
rect 95 -29 97 -25
rect 101 -29 103 -25
rect 105 -29 107 -25
rect 111 -29 113 -25
rect 115 -29 116 -25
rect 137 -29 138 -25
rect 140 -29 148 -25
rect 150 -29 152 -25
rect 156 -29 158 -25
rect 160 -29 161 -25
rect 181 -29 182 -25
rect 184 -29 192 -25
rect 194 -29 202 -25
rect 204 -29 205 -25
rect 214 -29 215 -25
rect 219 -29 220 -25
rect 222 -29 223 -25
rect 244 -29 245 -25
rect 247 -29 249 -25
rect 253 -29 255 -25
rect 257 -29 259 -25
rect 263 -29 265 -25
rect 267 -29 268 -25
rect 277 -29 278 -25
rect 282 -29 283 -25
rect 285 -29 286 -25
rect 309 -29 310 -25
rect 312 -29 320 -25
rect 322 -29 330 -25
rect 332 -29 341 -25
rect 343 -29 344 -25
rect 353 -29 354 -25
rect 358 -29 359 -25
rect 361 -29 362 -25
rect 384 -29 385 -25
rect 387 -29 395 -25
rect 397 -29 405 -25
rect 407 -29 408 -25
rect 417 -29 418 -25
rect 422 -29 423 -25
rect 425 -29 426 -25
rect 448 -29 449 -25
rect 451 -29 459 -25
rect 461 -29 463 -25
rect 467 -29 469 -25
rect 471 -29 472 -25
rect 493 -29 494 -25
rect 496 -29 498 -25
rect 502 -29 504 -25
rect 506 -29 508 -25
rect 512 -29 514 -25
rect 516 -29 519 -25
rect 523 -29 525 -25
rect 527 -29 528 -25
rect 537 -29 538 -25
rect 542 -29 543 -25
rect 545 -29 546 -25
<< pdiffusion >>
rect 42 4 43 12
rect 45 4 47 12
rect 51 4 53 12
rect 55 4 57 12
rect 61 4 63 12
rect 65 4 66 12
rect 92 4 93 12
rect 95 4 103 12
rect 105 4 107 12
rect 111 4 113 12
rect 115 4 116 12
rect 137 4 138 12
rect 140 4 142 12
rect 146 4 148 12
rect 150 4 152 12
rect 156 4 158 12
rect 160 4 161 12
rect 181 4 182 12
rect 184 4 186 12
rect 190 4 192 12
rect 194 4 196 12
rect 200 4 202 12
rect 204 4 205 12
rect 213 4 215 12
rect 219 4 220 12
rect 222 4 223 12
rect 244 4 245 12
rect 247 4 255 12
rect 257 4 265 12
rect 267 4 268 12
rect 277 4 278 12
rect 282 4 283 12
rect 285 4 286 12
rect 309 4 310 12
rect 312 4 314 12
rect 318 4 320 12
rect 322 4 324 12
rect 328 4 330 12
rect 332 4 334 12
rect 338 4 341 12
rect 343 4 344 12
rect 353 4 354 12
rect 358 4 359 12
rect 361 4 362 12
rect 384 4 385 12
rect 387 4 389 12
rect 393 4 395 12
rect 397 4 399 12
rect 403 4 405 12
rect 407 4 408 12
rect 416 4 418 12
rect 422 4 423 12
rect 425 4 426 12
rect 448 4 449 12
rect 451 4 453 12
rect 457 4 459 12
rect 461 4 463 12
rect 467 4 469 12
rect 471 4 472 12
rect 493 4 494 12
rect 496 4 504 12
rect 506 4 514 12
rect 516 4 525 12
rect 527 4 528 12
rect 537 4 538 12
rect 542 4 543 12
rect 545 4 546 12
<< ndcontact >>
rect 38 -29 42 -25
rect 57 -29 61 -25
rect 66 -29 70 -25
rect 88 -29 92 -25
rect 97 -29 101 -25
rect 107 -29 111 -25
rect 116 -29 120 -25
rect 133 -29 137 -25
rect 152 -29 156 -25
rect 161 -29 165 -25
rect 177 -29 181 -25
rect 205 -29 209 -25
rect 215 -29 219 -25
rect 223 -29 227 -25
rect 240 -29 244 -25
rect 249 -29 253 -25
rect 259 -29 263 -25
rect 268 -29 272 -25
rect 278 -29 282 -25
rect 286 -29 290 -25
rect 305 -29 309 -25
rect 344 -29 348 -25
rect 354 -29 358 -25
rect 362 -29 366 -25
rect 380 -29 384 -25
rect 408 -29 412 -25
rect 418 -29 422 -25
rect 426 -29 430 -25
rect 444 -29 448 -25
rect 463 -29 467 -25
rect 472 -29 476 -25
rect 489 -29 493 -25
rect 498 -29 502 -25
rect 508 -29 512 -25
rect 519 -29 523 -25
rect 528 -29 532 -25
rect 538 -29 542 -25
rect 546 -29 550 -25
<< pdcontact >>
rect 38 4 42 12
rect 47 4 51 12
rect 57 4 61 12
rect 66 4 70 12
rect 88 4 92 12
rect 107 4 111 12
rect 116 4 120 12
rect 133 4 137 12
rect 142 4 146 12
rect 152 4 156 12
rect 161 4 165 12
rect 177 4 181 12
rect 186 4 190 12
rect 196 4 200 12
rect 205 4 209 12
rect 215 4 219 12
rect 223 4 227 12
rect 240 4 244 12
rect 268 4 272 12
rect 278 4 282 12
rect 286 4 290 12
rect 305 4 309 12
rect 314 4 318 12
rect 324 4 328 12
rect 334 4 338 12
rect 344 4 348 12
rect 354 4 358 12
rect 362 4 366 12
rect 380 4 384 12
rect 389 4 393 12
rect 399 4 403 12
rect 408 4 412 12
rect 418 4 422 12
rect 426 4 430 12
rect 444 4 448 12
rect 453 4 457 12
rect 463 4 467 12
rect 472 4 476 12
rect 489 4 493 12
rect 528 4 532 12
rect 538 4 542 12
rect 546 4 550 12
<< psubstratepcontact >>
rect 37 -37 41 -33
rect 66 -37 70 -33
rect 87 -37 91 -33
rect 116 -37 120 -33
rect 132 -37 136 -33
rect 161 -37 165 -33
rect 176 -37 180 -33
rect 205 -37 209 -33
rect 227 -37 231 -33
rect 240 -37 244 -33
rect 268 -37 272 -33
rect 290 -37 294 -33
rect 305 -37 309 -33
rect 335 -37 339 -33
rect 366 -37 370 -33
rect 379 -37 383 -33
rect 408 -37 412 -33
rect 430 -37 434 -33
rect 443 -37 447 -33
rect 472 -37 476 -33
rect 489 -37 493 -33
rect 519 -37 523 -33
rect 550 -37 554 -33
<< nsubstratencontact >>
rect 38 17 42 21
rect 67 17 71 21
rect 88 17 92 21
rect 117 17 121 21
rect 133 17 137 21
rect 162 17 166 21
rect 177 17 181 21
rect 206 17 210 21
rect 225 17 229 21
rect 240 17 244 21
rect 269 17 273 21
rect 288 17 292 21
rect 305 17 309 21
rect 336 17 340 21
rect 364 17 368 21
rect 380 17 384 21
rect 409 17 413 21
rect 428 17 432 21
rect 444 17 448 21
rect 473 17 477 21
rect 489 17 493 21
rect 520 17 524 21
rect 548 17 552 21
<< polysilicon >>
rect 43 12 45 28
rect 53 12 55 28
rect 63 12 65 15
rect 93 12 95 15
rect 103 12 105 28
rect 113 12 115 15
rect 138 12 140 28
rect 148 12 150 28
rect 158 12 160 15
rect 182 12 184 28
rect 192 12 194 15
rect 202 12 204 28
rect 220 12 222 15
rect 245 12 247 15
rect 255 12 257 28
rect 265 12 267 15
rect 283 12 285 15
rect 310 12 312 15
rect 320 12 322 15
rect 330 12 332 28
rect 341 12 343 28
rect 359 12 361 15
rect 385 12 387 28
rect 395 12 397 15
rect 405 12 407 28
rect 423 12 425 15
rect 449 12 451 26
rect 459 12 461 26
rect 469 12 471 15
rect 494 12 496 15
rect 504 12 506 15
rect 514 12 516 15
rect 525 12 527 29
rect 543 12 545 15
rect 43 -25 45 4
rect 53 -25 55 4
rect 63 -25 65 4
rect 93 -25 95 4
rect 103 -25 105 4
rect 113 -25 115 4
rect 138 -25 140 4
rect 148 -25 150 4
rect 158 -25 160 4
rect 182 -25 184 4
rect 192 -25 194 4
rect 202 -25 204 4
rect 220 -25 222 4
rect 245 -25 247 4
rect 255 -25 257 4
rect 265 -25 267 4
rect 283 -25 285 4
rect 310 -25 312 4
rect 320 -25 322 4
rect 330 -25 332 4
rect 341 -25 343 4
rect 359 -25 361 4
rect 385 -25 387 4
rect 395 -25 397 4
rect 405 -25 407 4
rect 423 -25 425 4
rect 449 -25 451 4
rect 459 -25 461 4
rect 469 -25 471 4
rect 494 -25 496 4
rect 504 -25 506 4
rect 514 -25 516 4
rect 525 -25 527 4
rect 543 -25 545 4
rect 43 -32 45 -29
rect 53 -45 55 -29
rect 63 -32 65 -29
rect 93 -32 95 -29
rect 103 -32 105 -29
rect 113 -32 115 -29
rect 138 -32 140 -29
rect 148 -32 150 -29
rect 158 -32 160 -29
rect 182 -32 184 -29
rect 192 -46 194 -29
rect 202 -46 204 -29
rect 220 -32 222 -29
rect 245 -32 247 -29
rect 255 -32 257 -29
rect 265 -32 267 -29
rect 283 -32 285 -29
rect 310 -44 312 -29
rect 320 -44 322 -29
rect 330 -32 332 -29
rect 341 -32 343 -29
rect 359 -32 361 -29
rect 385 -32 387 -29
rect 395 -44 397 -29
rect 405 -32 407 -29
rect 423 -32 425 -29
rect 449 -32 451 -29
rect 459 -32 461 -29
rect 469 -32 471 -29
rect 494 -32 496 -29
rect 504 -32 506 -29
rect 514 -40 516 -29
rect 525 -32 527 -29
rect 543 -32 545 -29
<< polycontact >>
rect 39 24 43 28
rect 55 24 59 28
rect 105 24 109 28
rect 134 24 138 28
rect 150 24 154 28
rect 178 24 182 28
rect 204 24 208 28
rect 257 24 261 28
rect 332 24 336 28
rect 343 24 347 28
rect 381 24 385 28
rect 401 24 405 28
rect 448 26 452 30
rect 458 26 462 30
rect 521 24 525 28
rect 59 -8 63 -4
rect 89 -22 93 -18
rect 109 -16 113 -12
rect 154 -8 158 -4
rect 216 -19 220 -15
rect 241 -9 245 -5
rect 261 -9 265 -5
rect 279 -19 283 -15
rect 355 -19 359 -15
rect 419 -19 423 -15
rect 465 -8 469 -4
rect 490 -22 494 -18
rect 500 -9 504 -5
rect 539 -19 543 -15
rect 55 -44 59 -40
rect 188 -44 192 -40
rect 204 -44 208 -40
rect 306 -44 310 -40
rect 316 -44 320 -40
rect 391 -44 395 -40
rect 513 -44 517 -40
<< metal1 >>
rect -48 40 -43 47
rect 18 40 23 47
rect 18 28 23 35
rect 65 28 70 48
rect 117 47 120 48
rect 146 47 154 48
rect 146 44 208 47
rect 314 44 321 50
rect 362 46 366 50
rect 146 43 154 44
rect 116 28 121 42
rect 151 28 154 43
rect 179 28 182 34
rect 205 28 208 44
rect 317 31 320 44
rect 363 39 366 46
rect 467 47 472 52
rect 363 34 365 39
rect 18 24 39 28
rect 59 24 70 28
rect 109 24 134 28
rect 261 26 317 27
rect 333 28 336 34
rect 261 24 322 26
rect 363 27 366 34
rect 401 28 404 43
rect 347 24 381 27
rect 459 30 462 32
rect 442 27 448 30
rect 468 27 472 47
rect 468 24 521 27
rect 42 17 67 21
rect 71 17 88 21
rect 92 17 117 21
rect 121 17 133 21
rect 137 17 162 21
rect 166 17 177 21
rect 181 17 206 21
rect 210 17 225 21
rect 229 17 240 21
rect 244 17 269 21
rect 273 17 288 21
rect 292 17 305 21
rect 309 17 336 21
rect 340 17 364 21
rect 368 17 380 21
rect 384 17 409 21
rect 413 17 428 21
rect 432 17 444 21
rect 448 17 473 21
rect 477 17 489 21
rect 493 17 520 21
rect 524 17 548 21
rect 38 12 42 17
rect 57 12 61 17
rect 107 12 111 17
rect 133 12 137 17
rect 152 12 156 17
rect 177 12 181 17
rect 196 12 200 17
rect 215 12 219 17
rect 240 12 244 17
rect 278 12 282 17
rect 305 12 309 17
rect 324 12 328 17
rect 344 12 348 17
rect 47 -4 51 4
rect 47 -8 59 -4
rect 57 -18 61 -8
rect 38 -22 61 -18
rect 66 -19 70 4
rect 354 12 358 17
rect 380 12 384 17
rect 399 12 403 17
rect 418 12 422 17
rect 444 12 448 17
rect 463 12 467 17
rect 489 12 493 17
rect 538 12 542 17
rect 88 -12 92 4
rect 116 -8 120 4
rect 142 -4 146 4
rect 142 -8 154 -4
rect 88 -15 109 -12
rect 66 -22 89 -19
rect 38 -25 42 -22
rect 66 -25 70 -22
rect 97 -25 101 -15
rect 116 -13 121 -8
rect 116 -25 120 -13
rect 152 -18 156 -8
rect 133 -22 156 -18
rect 161 -17 165 4
rect 186 -4 190 4
rect 205 -4 209 4
rect 186 -8 209 -4
rect 205 -15 209 -8
rect 223 -13 227 4
rect 235 -9 241 -6
rect 259 -9 261 -5
rect 259 -13 262 -9
rect 161 -22 164 -17
rect 205 -19 216 -15
rect 223 -16 262 -13
rect 268 -15 272 4
rect 286 -9 290 4
rect 314 -8 318 4
rect 334 -8 338 4
rect 286 -13 292 -9
rect 314 -11 348 -8
rect 133 -25 137 -22
rect 161 -25 165 -22
rect 205 -25 209 -19
rect 223 -25 227 -16
rect 268 -19 279 -15
rect 249 -22 272 -19
rect 249 -25 253 -22
rect 268 -25 272 -22
rect 286 -25 290 -13
rect 344 -15 348 -11
rect 344 -19 355 -15
rect 344 -25 348 -19
rect 362 -25 366 4
rect 389 -4 393 4
rect 408 -4 412 4
rect 389 -8 412 -4
rect 408 -15 412 -8
rect 408 -19 419 -15
rect 426 -16 430 4
rect 453 -4 457 4
rect 453 -8 465 -4
rect 408 -25 412 -19
rect 426 -21 427 -16
rect 463 -18 467 -8
rect 426 -25 430 -21
rect 444 -22 467 -18
rect 472 -18 476 4
rect 491 -9 500 -6
rect 528 -15 532 4
rect 546 -9 550 4
rect 546 -13 552 -9
rect 472 -22 490 -18
rect 528 -19 539 -15
rect 498 -22 532 -19
rect 444 -25 448 -22
rect 472 -25 476 -22
rect 498 -25 502 -22
rect 519 -25 523 -22
rect 546 -25 550 -13
rect 57 -33 61 -29
rect 88 -33 92 -29
rect 107 -33 111 -29
rect 152 -33 156 -29
rect 177 -33 181 -29
rect 215 -33 219 -29
rect 240 -33 244 -29
rect 259 -33 263 -29
rect 278 -33 282 -29
rect 305 -33 309 -29
rect 354 -33 358 -29
rect 380 -33 384 -29
rect 418 -33 422 -29
rect 463 -33 467 -29
rect 489 -33 493 -29
rect 508 -33 512 -29
rect 528 -33 532 -29
rect 538 -33 542 -29
rect 41 -37 66 -33
rect 70 -37 87 -33
rect 91 -37 116 -33
rect 120 -37 132 -33
rect 136 -37 161 -33
rect 165 -37 176 -33
rect 180 -37 205 -33
rect 209 -37 227 -33
rect 231 -37 240 -33
rect 244 -37 268 -33
rect 272 -37 290 -33
rect 294 -37 305 -33
rect 309 -37 335 -33
rect 339 -37 366 -33
rect 370 -37 379 -33
rect 383 -37 408 -33
rect 412 -37 430 -33
rect 434 -37 443 -33
rect 447 -37 472 -33
rect 476 -37 489 -33
rect 493 -37 519 -33
rect 523 -37 550 -33
rect 59 -44 188 -41
rect 208 -41 306 -40
rect 208 -43 298 -41
rect 189 -49 192 -44
rect 303 -43 306 -41
rect 317 -49 320 -44
rect 388 -44 391 -41
rect 510 -44 513 -41
rect 189 -52 320 -49
<< m2contact >>
rect 18 35 23 40
rect 116 42 121 47
rect 179 34 184 39
rect 401 43 406 48
rect 332 34 337 39
rect 365 34 370 39
rect 317 26 322 31
rect 459 32 464 37
rect 437 27 442 32
rect 230 -9 235 -4
rect 164 -22 169 -17
rect 366 -10 371 -5
rect 427 -21 432 -16
rect 486 -10 491 -5
rect 298 -46 303 -41
rect 383 -45 388 -40
rect 505 -46 510 -41
<< metal2 >>
rect 19 44 23 49
rect 121 43 401 46
rect 23 35 179 38
rect 184 35 332 38
rect 370 37 463 39
rect 370 36 459 37
rect 322 27 437 30
rect 165 -9 230 -6
rect 165 -17 168 -9
rect 371 -10 486 -7
rect 303 -44 383 -41
rect 427 -41 430 -21
rect 427 -44 505 -41
<< labels >>
rlabel metal1 -47 47 -44 47 4 p0
rlabel m2contact 118 47 121 47 6 g1
rlabel metal1 121 -13 121 -8 1 c2
rlabel metal1 147 48 151 48 6 p2
rlabel metal1 255 19 255 19 5 vdd
rlabel metal1 256 -35 256 -35 1 gnd
rlabel metal1 292 -13 292 -9 1 c3
rlabel metal1 19 47 22 47 6 g0
rlabel metal1 316 50 320 50 6 g2
rlabel metal1 363 50 366 50 1 p3
rlabel metal1 468 52 472 52 1 g3
rlabel metal1 67 47 70 47 5 p1
rlabel metal1 552 -13 552 -9 1 c4
<< end >>
