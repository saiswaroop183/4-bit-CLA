magic
tech scmos
timestamp 1638596913
<< nwell >>
rect 32 -3 298 24
<< ntransistor >>
rect 43 -29 45 -25
rect 53 -29 55 -25
rect 63 -29 65 -25
rect 93 -29 95 -25
rect 103 -29 105 -25
rect 113 -29 115 -25
rect 138 -29 140 -25
rect 148 -29 150 -25
rect 158 -29 160 -25
rect 182 -29 184 -25
rect 192 -29 194 -25
rect 202 -29 204 -25
rect 220 -29 222 -25
rect 245 -29 247 -25
rect 255 -29 257 -25
rect 265 -29 267 -25
rect 283 -29 285 -25
<< ptransistor >>
rect 43 4 45 12
rect 53 4 55 12
rect 63 4 65 12
rect 93 4 95 12
rect 103 4 105 12
rect 113 4 115 12
rect 138 4 140 12
rect 148 4 150 12
rect 158 4 160 12
rect 182 4 184 12
rect 192 4 194 12
rect 202 4 204 12
rect 220 4 222 12
rect 245 4 247 12
rect 255 4 257 12
rect 265 4 267 12
rect 283 4 285 12
<< ndiffusion >>
rect 42 -29 43 -25
rect 45 -29 53 -25
rect 55 -29 57 -25
rect 61 -29 63 -25
rect 65 -29 66 -25
rect 92 -29 93 -25
rect 95 -29 97 -25
rect 101 -29 103 -25
rect 105 -29 107 -25
rect 111 -29 113 -25
rect 115 -29 116 -25
rect 137 -29 138 -25
rect 140 -29 148 -25
rect 150 -29 152 -25
rect 156 -29 158 -25
rect 160 -29 161 -25
rect 181 -29 182 -25
rect 184 -29 192 -25
rect 194 -29 202 -25
rect 204 -29 205 -25
rect 214 -29 215 -25
rect 219 -29 220 -25
rect 222 -29 223 -25
rect 244 -29 245 -25
rect 247 -29 249 -25
rect 253 -29 255 -25
rect 257 -29 259 -25
rect 263 -29 265 -25
rect 267 -29 268 -25
rect 277 -29 278 -25
rect 282 -29 283 -25
rect 285 -29 286 -25
<< pdiffusion >>
rect 42 4 43 12
rect 45 4 47 12
rect 51 4 53 12
rect 55 4 57 12
rect 61 4 63 12
rect 65 4 66 12
rect 92 4 93 12
rect 95 4 103 12
rect 105 4 107 12
rect 111 4 113 12
rect 115 4 116 12
rect 137 4 138 12
rect 140 4 142 12
rect 146 4 148 12
rect 150 4 152 12
rect 156 4 158 12
rect 160 4 161 12
rect 181 4 182 12
rect 184 4 186 12
rect 190 4 192 12
rect 194 4 196 12
rect 200 4 202 12
rect 204 4 205 12
rect 213 4 215 12
rect 219 4 220 12
rect 222 4 223 12
rect 244 4 245 12
rect 247 4 255 12
rect 257 4 265 12
rect 267 4 268 12
rect 277 4 278 12
rect 282 4 283 12
rect 285 4 286 12
<< ndcontact >>
rect 38 -29 42 -25
rect 57 -29 61 -25
rect 66 -29 70 -25
rect 88 -29 92 -25
rect 97 -29 101 -25
rect 107 -29 111 -25
rect 116 -29 120 -25
rect 133 -29 137 -25
rect 152 -29 156 -25
rect 161 -29 165 -25
rect 177 -29 181 -25
rect 205 -29 209 -25
rect 215 -29 219 -25
rect 223 -29 227 -25
rect 240 -29 244 -25
rect 249 -29 253 -25
rect 259 -29 263 -25
rect 268 -29 272 -25
rect 278 -29 282 -25
rect 286 -29 290 -25
<< pdcontact >>
rect 38 4 42 12
rect 47 4 51 12
rect 57 4 61 12
rect 66 4 70 12
rect 88 4 92 12
rect 107 4 111 12
rect 116 4 120 12
rect 133 4 137 12
rect 142 4 146 12
rect 152 4 156 12
rect 161 4 165 12
rect 177 4 181 12
rect 186 4 190 12
rect 196 4 200 12
rect 205 4 209 12
rect 215 4 219 12
rect 223 4 227 12
rect 240 4 244 12
rect 268 4 272 12
rect 278 4 282 12
rect 286 4 290 12
<< psubstratepcontact >>
rect 37 -37 41 -33
rect 66 -37 70 -33
rect 87 -37 91 -33
rect 116 -37 120 -33
rect 132 -37 136 -33
rect 161 -37 165 -33
rect 176 -37 180 -33
rect 205 -37 209 -33
rect 227 -37 231 -33
rect 240 -37 244 -33
rect 268 -37 272 -33
rect 290 -37 294 -33
<< nsubstratencontact >>
rect 38 17 42 21
rect 67 17 71 21
rect 88 17 92 21
rect 117 17 121 21
rect 133 17 137 21
rect 162 17 166 21
rect 177 17 181 21
rect 206 17 210 21
rect 225 17 229 21
rect 240 17 244 21
rect 269 17 273 21
rect 288 17 292 21
<< polysilicon >>
rect 43 12 45 28
rect 53 12 55 28
rect 63 12 65 15
rect 93 12 95 15
rect 103 12 105 28
rect 113 12 115 15
rect 138 12 140 28
rect 148 12 150 28
rect 158 12 160 15
rect 182 12 184 28
rect 192 12 194 15
rect 202 12 204 28
rect 220 12 222 15
rect 245 12 247 15
rect 255 12 257 28
rect 265 12 267 15
rect 283 12 285 15
rect 43 -25 45 4
rect 53 -25 55 4
rect 63 -25 65 4
rect 93 -25 95 4
rect 103 -25 105 4
rect 113 -25 115 4
rect 138 -25 140 4
rect 148 -25 150 4
rect 158 -25 160 4
rect 182 -25 184 4
rect 192 -25 194 4
rect 202 -25 204 4
rect 220 -25 222 4
rect 245 -25 247 4
rect 255 -25 257 4
rect 265 -25 267 4
rect 283 -25 285 4
rect 43 -32 45 -29
rect 53 -45 55 -29
rect 63 -32 65 -29
rect 93 -32 95 -29
rect 103 -32 105 -29
rect 113 -32 115 -29
rect 138 -32 140 -29
rect 148 -32 150 -29
rect 158 -32 160 -29
rect 182 -32 184 -29
rect 192 -46 194 -29
rect 202 -32 204 -29
rect 220 -32 222 -29
rect 245 -32 247 -29
rect 255 -32 257 -29
rect 265 -32 267 -29
rect 283 -32 285 -29
<< polycontact >>
rect 39 24 43 28
rect 55 24 59 28
rect 105 24 109 28
rect 134 24 138 28
rect 150 24 154 28
rect 178 24 182 28
rect 204 24 208 28
rect 251 24 255 28
rect 59 -8 63 -4
rect 89 -22 93 -18
rect 109 -16 113 -12
rect 154 -8 158 -4
rect 216 -19 220 -15
rect 241 -9 245 -5
rect 261 -9 265 -5
rect 279 -19 283 -15
rect 55 -44 59 -40
rect 188 -44 192 -40
<< metal1 >>
rect 146 47 154 48
rect -48 40 -43 47
rect 18 44 23 47
rect 18 28 23 39
rect 65 28 70 47
rect 116 28 121 47
rect 146 44 208 47
rect 146 43 154 44
rect 151 28 154 43
rect 179 28 182 34
rect 205 28 208 44
rect 219 42 226 48
rect 18 24 39 28
rect 59 24 70 28
rect 109 24 134 28
rect 222 27 225 42
rect 222 24 251 27
rect 42 17 67 21
rect 71 17 88 21
rect 92 17 117 21
rect 121 17 133 21
rect 137 17 162 21
rect 166 17 177 21
rect 181 17 206 21
rect 210 17 225 21
rect 229 17 240 21
rect 244 17 269 21
rect 273 17 288 21
rect 38 12 42 17
rect 57 12 61 17
rect 107 12 111 17
rect 133 12 137 17
rect 152 12 156 17
rect 177 12 181 17
rect 196 12 200 17
rect 215 12 219 17
rect 240 12 244 17
rect 278 12 282 17
rect 47 -4 51 4
rect 47 -8 59 -4
rect 57 -18 61 -8
rect 38 -22 61 -18
rect 66 -19 70 4
rect 88 -12 92 4
rect 116 -8 120 4
rect 142 -4 146 4
rect 142 -8 154 -4
rect 88 -15 109 -12
rect 66 -22 89 -19
rect 38 -25 42 -22
rect 66 -25 70 -22
rect 97 -25 101 -15
rect 116 -13 121 -8
rect 116 -25 120 -13
rect 152 -18 156 -8
rect 133 -22 156 -18
rect 161 -17 165 4
rect 186 -4 190 4
rect 205 -4 209 4
rect 186 -8 209 -4
rect 205 -15 209 -8
rect 223 -13 227 4
rect 235 -9 241 -6
rect 259 -9 261 -5
rect 259 -13 262 -9
rect 161 -22 164 -17
rect 205 -19 216 -15
rect 223 -16 262 -13
rect 268 -15 272 4
rect 286 -9 290 4
rect 286 -13 292 -9
rect 133 -25 137 -22
rect 161 -25 165 -22
rect 205 -25 209 -19
rect 223 -25 227 -16
rect 268 -19 279 -15
rect 249 -22 272 -19
rect 249 -25 253 -22
rect 268 -25 272 -22
rect 286 -25 290 -13
rect 57 -33 61 -29
rect 88 -33 92 -29
rect 107 -33 111 -29
rect 152 -33 156 -29
rect 177 -33 181 -29
rect 215 -33 219 -29
rect 240 -33 244 -29
rect 259 -33 263 -29
rect 278 -33 282 -29
rect 41 -37 66 -33
rect 70 -37 87 -33
rect 91 -37 116 -33
rect 120 -37 132 -33
rect 136 -37 161 -33
rect 165 -37 176 -33
rect 180 -37 205 -33
rect 209 -37 227 -33
rect 231 -37 240 -33
rect 244 -37 268 -33
rect 272 -37 290 -33
rect 59 -44 188 -41
<< m2contact >>
rect 18 39 23 44
rect 179 34 184 39
rect 230 -9 235 -4
rect 164 -22 169 -17
<< metal2 >>
rect 23 39 182 42
rect 165 -9 230 -6
rect 165 -17 168 -9
<< labels >>
rlabel metal1 -47 47 -44 47 4 p0
rlabel metal1 19 47 22 47 6 g0
rlabel metal1 67 47 70 47 5 p1
rlabel metal1 118 47 121 47 6 g1
rlabel metal1 121 -13 121 -8 1 c2
rlabel metal1 147 48 151 48 6 p2
rlabel metal1 221 48 225 48 6 g2
rlabel metal1 255 19 255 19 5 vdd
rlabel metal1 256 -35 256 -35 1 gnd
rlabel metal1 292 -13 292 -9 1 c3
<< end >>
