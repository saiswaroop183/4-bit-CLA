magic
tech scmos
timestamp 1638560381
<< nwell >>
rect -58 0 538 27
<< ntransistor >>
rect -47 -43 -45 -39
rect -34 -43 -32 -39
rect -16 -43 -14 -39
rect -6 -43 -4 -39
rect 13 -43 15 -39
rect 33 -43 35 -39
rect 102 -43 104 -39
rect 115 -43 117 -39
rect 133 -43 135 -39
rect 143 -43 145 -39
rect 162 -43 164 -39
rect 182 -43 184 -39
rect 251 -43 253 -39
rect 264 -43 266 -39
rect 282 -43 284 -39
rect 292 -43 294 -39
rect 311 -43 313 -39
rect 331 -43 333 -39
rect 400 -43 402 -39
rect 413 -43 415 -39
rect 431 -43 433 -39
rect 441 -43 443 -39
rect 460 -43 462 -39
rect 480 -43 482 -39
rect 57 -50 59 -46
rect 67 -50 69 -46
rect 77 -50 79 -46
rect 206 -50 208 -46
rect 216 -50 218 -46
rect 226 -50 228 -46
rect 355 -50 357 -46
rect 365 -50 367 -46
rect 375 -50 377 -46
rect 504 -50 506 -46
rect 514 -50 516 -46
rect 524 -50 526 -46
<< ptransistor >>
rect -47 7 -45 15
rect -34 7 -32 15
rect -16 7 -14 15
rect -6 7 -4 15
rect 13 7 15 15
rect 33 7 35 15
rect 57 7 59 15
rect 67 7 69 15
rect 77 7 79 15
rect 102 7 104 15
rect 115 7 117 15
rect 133 7 135 15
rect 143 7 145 15
rect 162 7 164 15
rect 182 7 184 15
rect 206 7 208 15
rect 216 7 218 15
rect 226 7 228 15
rect 251 7 253 15
rect 264 7 266 15
rect 282 7 284 15
rect 292 7 294 15
rect 311 7 313 15
rect 331 7 333 15
rect 355 7 357 15
rect 365 7 367 15
rect 375 7 377 15
rect 400 7 402 15
rect 413 7 415 15
rect 431 7 433 15
rect 441 7 443 15
rect 460 7 462 15
rect 480 7 482 15
rect 504 7 506 15
rect 514 7 516 15
rect 524 7 526 15
<< ndiffusion >>
rect -48 -43 -47 -39
rect -45 -43 -42 -39
rect -38 -43 -34 -39
rect -32 -43 -31 -39
rect -17 -43 -16 -39
rect -14 -43 -12 -39
rect -8 -43 -6 -39
rect -4 -43 -2 -39
rect 2 -43 13 -39
rect 15 -43 17 -39
rect 21 -43 33 -39
rect 35 -43 36 -39
rect 101 -43 102 -39
rect 104 -43 107 -39
rect 111 -43 115 -39
rect 117 -43 118 -39
rect 132 -43 133 -39
rect 135 -43 137 -39
rect 141 -43 143 -39
rect 145 -43 147 -39
rect 151 -43 162 -39
rect 164 -43 166 -39
rect 170 -43 182 -39
rect 184 -43 185 -39
rect 250 -43 251 -39
rect 253 -43 256 -39
rect 260 -43 264 -39
rect 266 -43 267 -39
rect 281 -43 282 -39
rect 284 -43 286 -39
rect 290 -43 292 -39
rect 294 -43 296 -39
rect 300 -43 311 -39
rect 313 -43 315 -39
rect 319 -43 331 -39
rect 333 -43 334 -39
rect 399 -43 400 -39
rect 402 -43 405 -39
rect 409 -43 413 -39
rect 415 -43 416 -39
rect 430 -43 431 -39
rect 433 -43 435 -39
rect 439 -43 441 -39
rect 443 -43 445 -39
rect 449 -43 460 -39
rect 462 -43 464 -39
rect 468 -43 480 -39
rect 482 -43 483 -39
rect 56 -50 57 -46
rect 59 -50 67 -46
rect 69 -50 71 -46
rect 75 -50 77 -46
rect 79 -50 80 -46
rect 205 -50 206 -46
rect 208 -50 216 -46
rect 218 -50 220 -46
rect 224 -50 226 -46
rect 228 -50 229 -46
rect 354 -50 355 -46
rect 357 -50 365 -46
rect 367 -50 369 -46
rect 373 -50 375 -46
rect 377 -50 378 -46
rect 503 -50 504 -46
rect 506 -50 514 -46
rect 516 -50 518 -46
rect 522 -50 524 -46
rect 526 -50 527 -46
<< pdiffusion >>
rect -48 7 -47 15
rect -45 7 -39 15
rect -35 7 -34 15
rect -32 7 -31 15
rect -17 7 -16 15
rect -14 7 -6 15
rect -4 7 -2 15
rect 2 7 13 15
rect 15 7 33 15
rect 35 7 36 15
rect 56 7 57 15
rect 59 7 61 15
rect 65 7 67 15
rect 69 7 71 15
rect 75 7 77 15
rect 79 7 80 15
rect 101 7 102 15
rect 104 7 110 15
rect 114 7 115 15
rect 117 7 118 15
rect 132 7 133 15
rect 135 7 143 15
rect 145 7 147 15
rect 151 7 162 15
rect 164 7 182 15
rect 184 7 185 15
rect 205 7 206 15
rect 208 7 210 15
rect 214 7 216 15
rect 218 7 220 15
rect 224 7 226 15
rect 228 7 229 15
rect 250 7 251 15
rect 253 7 259 15
rect 263 7 264 15
rect 266 7 267 15
rect 281 7 282 15
rect 284 7 292 15
rect 294 7 296 15
rect 300 7 311 15
rect 313 7 331 15
rect 333 7 334 15
rect 354 7 355 15
rect 357 7 359 15
rect 363 7 365 15
rect 367 7 369 15
rect 373 7 375 15
rect 377 7 378 15
rect 399 7 400 15
rect 402 7 408 15
rect 412 7 413 15
rect 415 7 416 15
rect 430 7 431 15
rect 433 7 441 15
rect 443 7 445 15
rect 449 7 460 15
rect 462 7 480 15
rect 482 7 483 15
rect 503 7 504 15
rect 506 7 508 15
rect 512 7 514 15
rect 516 7 518 15
rect 522 7 524 15
rect 526 7 527 15
<< ndcontact >>
rect -52 -43 -48 -39
rect -42 -43 -38 -39
rect -31 -43 -27 -39
rect -21 -43 -17 -39
rect -12 -43 -8 -39
rect -2 -43 2 -39
rect 17 -43 21 -39
rect 36 -43 40 -39
rect 97 -43 101 -39
rect 107 -43 111 -39
rect 118 -43 122 -39
rect 128 -43 132 -39
rect 137 -43 141 -39
rect 147 -43 151 -39
rect 166 -43 170 -39
rect 185 -43 189 -39
rect 246 -43 250 -39
rect 256 -43 260 -39
rect 267 -43 271 -39
rect 277 -43 281 -39
rect 286 -43 290 -39
rect 296 -43 300 -39
rect 315 -43 319 -39
rect 334 -43 338 -39
rect 395 -43 399 -39
rect 405 -43 409 -39
rect 416 -43 420 -39
rect 426 -43 430 -39
rect 435 -43 439 -39
rect 445 -43 449 -39
rect 464 -43 468 -39
rect 483 -43 487 -39
rect 52 -50 56 -46
rect 71 -50 75 -46
rect 80 -50 84 -46
rect 201 -50 205 -46
rect 220 -50 224 -46
rect 229 -50 233 -46
rect 350 -50 354 -46
rect 369 -50 373 -46
rect 378 -50 382 -46
rect 499 -50 503 -46
rect 518 -50 522 -46
rect 527 -50 531 -46
<< pdcontact >>
rect -52 7 -48 15
rect -39 7 -35 15
rect -31 7 -27 15
rect -21 7 -17 15
rect -2 7 2 15
rect 36 7 40 15
rect 52 7 56 15
rect 61 7 65 15
rect 71 7 75 15
rect 80 7 84 15
rect 97 7 101 15
rect 110 7 114 15
rect 118 7 122 15
rect 128 7 132 15
rect 147 7 151 15
rect 185 7 189 15
rect 201 7 205 15
rect 210 7 214 15
rect 220 7 224 15
rect 229 7 233 15
rect 246 7 250 15
rect 259 7 263 15
rect 267 7 271 15
rect 277 7 281 15
rect 296 7 300 15
rect 334 7 338 15
rect 350 7 354 15
rect 359 7 363 15
rect 369 7 373 15
rect 378 7 382 15
rect 395 7 399 15
rect 408 7 412 15
rect 416 7 420 15
rect 426 7 430 15
rect 445 7 449 15
rect 483 7 487 15
rect 499 7 503 15
rect 508 7 512 15
rect 518 7 522 15
rect 527 7 531 15
<< psubstratepcontact >>
rect -58 -58 -54 -54
rect -40 -58 -36 -54
rect -22 -58 -18 -54
rect 11 -58 15 -54
rect 41 -58 45 -54
rect 51 -58 55 -54
rect 80 -58 84 -54
rect 91 -58 95 -54
rect 109 -58 113 -54
rect 127 -58 131 -54
rect 160 -58 164 -54
rect 190 -58 194 -54
rect 200 -58 204 -54
rect 229 -58 233 -54
rect 240 -58 244 -54
rect 258 -58 262 -54
rect 276 -58 280 -54
rect 309 -58 313 -54
rect 339 -58 343 -54
rect 349 -58 353 -54
rect 378 -58 382 -54
rect 389 -58 393 -54
rect 407 -58 411 -54
rect 425 -58 429 -54
rect 458 -58 462 -54
rect 488 -58 492 -54
rect 498 -58 502 -54
rect 527 -58 531 -54
<< nsubstratencontact >>
rect -54 20 -50 24
rect -29 20 -25 24
rect -21 20 -17 24
rect -2 20 2 24
rect 39 20 43 24
rect 52 20 56 24
rect 81 20 85 24
rect 95 20 99 24
rect 120 20 124 24
rect 128 20 132 24
rect 147 20 151 24
rect 188 20 192 24
rect 201 20 205 24
rect 230 20 234 24
rect 244 20 248 24
rect 269 20 273 24
rect 277 20 281 24
rect 296 20 300 24
rect 337 20 341 24
rect 350 20 354 24
rect 379 20 383 24
rect 393 20 397 24
rect 418 20 422 24
rect 426 20 430 24
rect 445 20 449 24
rect 486 20 490 24
rect 499 20 503 24
rect 528 20 532 24
<< polysilicon >>
rect -47 15 -45 19
rect -34 15 -32 19
rect -16 15 -14 18
rect -6 15 -4 18
rect 13 15 15 18
rect 33 15 35 18
rect 57 15 59 18
rect 67 15 69 18
rect 77 15 79 18
rect 102 15 104 19
rect 115 15 117 19
rect 133 15 135 18
rect 143 15 145 18
rect 162 15 164 18
rect 182 15 184 18
rect 206 15 208 18
rect 216 15 218 18
rect 226 15 228 18
rect 251 15 253 19
rect 264 15 266 19
rect 282 15 284 18
rect 292 15 294 18
rect 311 15 313 18
rect 331 15 333 18
rect 355 15 357 18
rect 365 15 367 18
rect 375 15 377 18
rect 400 15 402 19
rect 413 15 415 19
rect 431 15 433 18
rect 441 15 443 18
rect 460 15 462 18
rect 480 15 482 18
rect 504 15 506 18
rect 514 15 516 18
rect 524 15 526 18
rect -47 -39 -45 7
rect -34 -39 -32 7
rect -16 -39 -14 7
rect -6 -39 -4 7
rect 13 -39 15 7
rect 33 -39 35 7
rect -47 -46 -45 -43
rect -34 -46 -32 -43
rect -16 -46 -14 -43
rect -6 -46 -4 -43
rect 13 -46 15 -43
rect 33 -46 35 -43
rect 57 -46 59 7
rect 67 -46 69 7
rect 77 -46 79 7
rect 102 -39 104 7
rect 115 -39 117 7
rect 133 -39 135 7
rect 143 -39 145 7
rect 162 -39 164 7
rect 182 -39 184 7
rect 102 -46 104 -43
rect 115 -46 117 -43
rect 133 -46 135 -43
rect 143 -46 145 -43
rect 162 -46 164 -43
rect 182 -46 184 -43
rect 206 -46 208 7
rect 216 -46 218 7
rect 226 -46 228 7
rect 251 -39 253 7
rect 264 -39 266 7
rect 282 -39 284 7
rect 292 -39 294 7
rect 311 -39 313 7
rect 331 -39 333 7
rect 251 -46 253 -43
rect 264 -46 266 -43
rect 282 -46 284 -43
rect 292 -46 294 -43
rect 311 -46 313 -43
rect 331 -46 333 -43
rect 355 -46 357 7
rect 365 -46 367 7
rect 375 -46 377 7
rect 400 -39 402 7
rect 413 -39 415 7
rect 431 -39 433 7
rect 441 -39 443 7
rect 460 -39 462 7
rect 480 -39 482 7
rect 400 -46 402 -43
rect 413 -46 415 -43
rect 431 -46 433 -43
rect 441 -46 443 -43
rect 460 -46 462 -43
rect 480 -46 482 -43
rect 504 -46 506 7
rect 514 -46 516 7
rect 524 -46 526 7
rect 57 -53 59 -50
rect 67 -53 69 -50
rect 77 -53 79 -50
rect 206 -53 208 -50
rect 216 -53 218 -50
rect 226 -53 228 -50
rect 355 -53 357 -50
rect 365 -53 367 -50
rect 375 -53 377 -50
rect 504 -53 506 -50
rect 514 -53 516 -50
rect 524 -53 526 -50
<< polycontact >>
rect -45 -9 -41 -5
rect -38 -35 -34 -31
rect -20 -34 -16 -30
rect -4 -16 0 -12
rect 15 -18 19 -14
rect 53 -6 57 -2
rect 35 -22 39 -18
rect 63 -12 67 -8
rect 73 -5 77 -1
rect 104 -9 108 -5
rect 111 -35 115 -31
rect 129 -34 133 -30
rect 145 -16 149 -12
rect 164 -18 168 -14
rect 202 -6 206 -2
rect 184 -22 188 -18
rect 212 -12 216 -8
rect 222 -5 226 -1
rect 253 -9 257 -5
rect 260 -35 264 -31
rect 278 -34 282 -30
rect 294 -16 298 -12
rect 313 -18 317 -14
rect 351 -6 355 -2
rect 333 -22 337 -18
rect 361 -12 365 -8
rect 371 -5 375 -1
rect 402 -9 406 -5
rect 409 -35 413 -31
rect 427 -34 431 -30
rect 443 -16 447 -12
rect 462 -18 466 -14
rect 500 -6 504 -2
rect 482 -22 486 -18
rect 510 -12 514 -8
rect 520 -5 524 -1
<< metal1 >>
rect -50 20 -29 24
rect -25 20 -21 24
rect -17 20 -2 24
rect 2 20 39 24
rect 43 20 52 24
rect 56 20 81 24
rect 85 20 95 24
rect 99 20 120 24
rect 124 20 128 24
rect 132 20 147 24
rect 151 20 188 24
rect 192 20 201 24
rect 205 20 230 24
rect 234 20 244 24
rect 248 20 269 24
rect 273 20 277 24
rect 281 20 296 24
rect 300 20 337 24
rect 341 20 350 24
rect 354 20 379 24
rect 383 20 393 24
rect 397 20 418 24
rect 422 20 426 24
rect 430 20 445 24
rect 449 20 486 24
rect 490 20 499 24
rect 503 20 528 24
rect -39 15 -35 20
rect -2 15 2 20
rect 52 15 56 20
rect 71 15 75 20
rect 110 15 114 20
rect 147 15 151 20
rect 201 15 205 20
rect 220 15 224 20
rect 259 15 263 20
rect 296 15 300 20
rect 350 15 354 20
rect 369 15 373 20
rect 408 15 412 20
rect 445 15 449 20
rect 499 15 503 20
rect 518 15 522 20
rect -52 -33 -48 7
rect -41 -9 -40 -5
rect -31 -30 -27 7
rect -21 -2 -17 7
rect 36 -2 40 7
rect 61 -1 65 7
rect -21 -7 40 -2
rect 48 -3 53 -2
rect -12 -11 -8 -7
rect 49 -7 53 -3
rect 61 -5 73 -1
rect 0 -16 1 -12
rect -55 -37 -48 -33
rect -39 -35 -38 -31
rect -31 -34 -20 -30
rect -52 -39 -48 -37
rect -31 -39 -27 -34
rect -12 -39 -8 -16
rect 19 -18 23 -14
rect 60 -18 63 -8
rect 39 -22 43 -18
rect 48 -22 63 -18
rect -2 -36 40 -32
rect -2 -39 2 -36
rect 36 -39 40 -36
rect 71 -39 75 -5
rect -42 -54 -38 -43
rect -21 -47 -17 -43
rect -2 -47 2 -43
rect -21 -51 2 -47
rect 52 -43 75 -39
rect 80 -9 84 7
rect 80 -13 86 -9
rect 17 -54 21 -43
rect 52 -46 56 -43
rect 80 -46 84 -13
rect 97 -33 101 7
rect 108 -9 109 -5
rect 118 -30 122 7
rect 128 -2 132 7
rect 185 -2 189 7
rect 210 -1 214 7
rect 128 -7 189 -2
rect 197 -3 202 -2
rect 137 -11 141 -7
rect 198 -7 202 -3
rect 210 -5 222 -1
rect 149 -16 150 -12
rect 94 -37 101 -33
rect 110 -35 111 -31
rect 118 -34 129 -30
rect 97 -39 101 -37
rect 118 -39 122 -34
rect 137 -39 141 -16
rect 168 -18 172 -14
rect 209 -18 212 -8
rect 188 -22 192 -18
rect 197 -22 212 -18
rect 147 -36 189 -32
rect 147 -39 151 -36
rect 185 -39 189 -36
rect 220 -39 224 -5
rect 71 -54 75 -50
rect 107 -54 111 -43
rect 128 -47 132 -43
rect 147 -47 151 -43
rect 128 -51 151 -47
rect 201 -43 224 -39
rect 229 -10 233 7
rect 229 -13 235 -10
rect 166 -54 170 -43
rect 201 -46 205 -43
rect 229 -46 233 -13
rect 246 -33 250 7
rect 257 -9 258 -5
rect 267 -30 271 7
rect 277 -2 281 7
rect 334 -2 338 7
rect 359 -1 363 7
rect 277 -7 338 -2
rect 346 -3 351 -2
rect 286 -11 290 -7
rect 347 -7 351 -3
rect 359 -5 371 -1
rect 298 -16 299 -12
rect 243 -37 250 -33
rect 259 -35 260 -31
rect 267 -34 278 -30
rect 246 -39 250 -37
rect 267 -39 271 -34
rect 286 -39 290 -16
rect 317 -18 321 -14
rect 358 -18 361 -8
rect 337 -22 341 -18
rect 346 -22 361 -18
rect 296 -36 338 -32
rect 296 -39 300 -36
rect 334 -39 338 -36
rect 369 -39 373 -5
rect 220 -54 224 -50
rect 256 -54 260 -43
rect 277 -47 281 -43
rect 296 -47 300 -43
rect 277 -51 300 -47
rect 350 -43 373 -39
rect 378 -10 382 7
rect 378 -13 384 -10
rect 315 -54 319 -43
rect 350 -46 354 -43
rect 378 -46 382 -13
rect 395 -33 399 7
rect 406 -9 407 -5
rect 416 -30 420 7
rect 426 -2 430 7
rect 483 -2 487 7
rect 508 -1 512 7
rect 426 -7 487 -2
rect 495 -3 500 -2
rect 435 -11 439 -7
rect 496 -7 500 -3
rect 508 -5 520 -1
rect 447 -16 448 -12
rect 392 -37 399 -33
rect 408 -35 409 -31
rect 416 -34 427 -30
rect 395 -39 399 -37
rect 416 -39 420 -34
rect 435 -39 439 -16
rect 466 -18 470 -14
rect 507 -18 510 -8
rect 486 -22 490 -18
rect 495 -22 510 -18
rect 445 -36 487 -32
rect 445 -39 449 -36
rect 483 -39 487 -36
rect 518 -39 522 -5
rect 369 -54 373 -50
rect 405 -54 409 -43
rect 426 -47 430 -43
rect 445 -47 449 -43
rect 426 -51 449 -47
rect 499 -43 522 -39
rect 527 -10 531 7
rect 527 -13 533 -10
rect 464 -54 468 -43
rect 499 -46 503 -43
rect 527 -46 531 -13
rect 518 -54 522 -50
rect -54 -58 -40 -54
rect -36 -58 -22 -54
rect -18 -58 11 -54
rect 15 -58 41 -54
rect 45 -58 51 -54
rect 55 -58 80 -54
rect 84 -58 91 -54
rect 95 -58 109 -54
rect 113 -58 127 -54
rect 131 -58 160 -54
rect 164 -58 190 -54
rect 194 -58 200 -54
rect 204 -58 229 -54
rect 233 -58 240 -54
rect 244 -58 258 -54
rect 262 -58 276 -54
rect 280 -58 309 -54
rect 313 -58 339 -54
rect 343 -58 349 -54
rect 353 -58 378 -54
rect 382 -58 389 -54
rect 393 -58 407 -54
rect 411 -58 425 -54
rect 429 -58 458 -54
rect 462 -58 488 -54
rect 492 -58 498 -54
rect 502 -58 527 -54
<< m2contact >>
rect -60 -37 -55 -32
rect -40 -9 -35 -4
rect 44 -8 49 -3
rect -12 -16 -7 -11
rect 1 -16 6 -11
rect -44 -35 -39 -30
rect 23 -19 28 -14
rect 43 -23 48 -18
rect 89 -37 94 -32
rect 109 -9 114 -4
rect 193 -8 198 -3
rect 137 -16 142 -11
rect 150 -16 155 -11
rect 105 -35 110 -30
rect 172 -19 177 -14
rect 192 -23 197 -18
rect 238 -37 243 -32
rect 258 -9 263 -4
rect 342 -8 347 -3
rect 286 -16 291 -11
rect 299 -16 304 -11
rect 254 -35 259 -30
rect 321 -19 326 -14
rect 341 -23 346 -18
rect 387 -37 392 -32
rect 407 -9 412 -4
rect 491 -8 496 -3
rect 435 -16 440 -11
rect 448 -16 453 -11
rect 403 -35 408 -30
rect 470 -19 475 -14
rect 490 -23 495 -18
<< metal2 >>
rect -62 -7 -40 -4
rect -35 -7 44 -4
rect 4 -8 44 -7
rect 87 -7 109 -4
rect 4 -11 8 -8
rect 114 -7 193 -4
rect 153 -8 193 -7
rect 236 -7 258 -4
rect 153 -11 157 -8
rect 263 -7 342 -4
rect 302 -8 342 -7
rect 385 -7 407 -4
rect 302 -11 306 -8
rect 412 -7 491 -4
rect 451 -8 491 -7
rect 451 -11 455 -8
rect -62 -16 -12 -13
rect 6 -16 8 -11
rect 87 -16 137 -13
rect 155 -16 157 -11
rect 23 -20 27 -19
rect -59 -23 27 -20
rect 236 -16 286 -13
rect 304 -16 306 -11
rect 172 -20 176 -19
rect 90 -23 176 -20
rect 385 -16 435 -13
rect 453 -16 455 -11
rect 321 -20 325 -19
rect 239 -23 325 -20
rect 470 -20 474 -19
rect 388 -23 474 -20
rect -59 -32 -56 -23
rect 43 -32 46 -23
rect 90 -32 93 -23
rect -39 -35 46 -32
rect -35 -47 -32 -35
rect 192 -32 195 -23
rect 239 -32 242 -23
rect 110 -35 195 -32
rect 114 -47 117 -35
rect 341 -32 344 -23
rect 388 -32 391 -23
rect 259 -35 344 -32
rect 263 -47 266 -35
rect 490 -32 493 -23
rect 408 -35 493 -32
rect 412 -47 415 -35
rect -62 -50 -32 -47
rect 87 -50 117 -47
rect 236 -50 266 -47
rect 385 -50 415 -47
<< labels >>
rlabel metal2 -61 -50 -61 -47 3 a0
rlabel metal1 86 -13 86 -9 7 g0
rlabel metal2 -62 -7 -62 -4 3 b0
rlabel metal2 -61 -16 -61 -13 3 p0
rlabel metal1 166 22 166 22 5 vdd
rlabel metal1 146 -56 146 -56 1 gnd
rlabel metal2 87 -7 87 -4 1 b1
rlabel metal2 88 -50 88 -47 1 a1
rlabel metal2 88 -16 88 -13 1 p1
rlabel metal1 235 -13 235 -10 1 g1
rlabel metal2 236 -7 236 -4 1 b2
rlabel metal2 237 -16 237 -13 1 p2
rlabel metal2 237 -50 237 -47 1 a2
rlabel metal1 384 -13 384 -10 1 g2
rlabel metal2 385 -7 385 -4 1 b3
rlabel metal2 386 -16 386 -13 1 p3
rlabel metal2 386 -50 386 -47 1 a3
rlabel metal1 533 -13 533 -10 7 g3
<< end >>
