magic
tech scmos
timestamp 1637319880
<< nwell >>
rect -27 0 18 27
<< ntransistor >>
rect -16 -20 -14 -16
rect -6 -20 -4 -16
rect 4 -20 6 -16
<< ptransistor >>
rect -16 7 -14 15
rect -6 7 -4 15
rect 4 7 6 15
<< ndiffusion >>
rect -17 -20 -16 -16
rect -14 -20 -12 -16
rect -8 -20 -6 -16
rect -4 -20 -2 -16
rect 2 -20 4 -16
rect 6 -20 7 -16
<< pdiffusion >>
rect -17 7 -16 15
rect -14 7 -6 15
rect -4 7 -2 15
rect 2 7 4 15
rect 6 7 7 15
<< ndcontact >>
rect -21 -20 -17 -16
rect -12 -20 -8 -16
rect -2 -20 2 -16
rect 7 -20 11 -16
<< pdcontact >>
rect -21 7 -17 15
rect -2 7 2 15
rect 7 7 11 15
<< psubstratepcontact >>
rect -22 -28 -18 -24
rect 7 -28 11 -24
<< nsubstratencontact >>
rect -21 20 -17 24
rect 8 20 12 24
<< polysilicon >>
rect -16 15 -14 18
rect -6 15 -4 18
rect 4 15 6 18
rect -16 -16 -14 7
rect -6 -16 -4 7
rect 4 -16 6 7
rect -16 -23 -14 -20
rect -6 -23 -4 -20
rect 4 -23 6 -20
<< polycontact >>
rect -14 -5 -10 -1
rect -4 -5 0 -1
rect 0 -13 4 -9
<< metal1 >>
rect -17 20 8 24
rect -2 15 2 20
rect -21 -9 -17 7
rect -10 -5 -8 -1
rect 0 -5 2 -1
rect 7 -5 11 7
rect -21 -13 0 -9
rect 7 -10 12 -5
rect -12 -16 -8 -13
rect 7 -16 11 -10
rect -21 -24 -17 -20
rect -2 -24 2 -20
rect -18 -28 7 -24
<< labels >>
rlabel metal1 12 -10 12 -5 1 g
rlabel metal1 -5 -26 -5 -26 1 gnd
rlabel metal1 -8 -5 -8 -1 1 a
rlabel metal1 2 -5 2 -1 1 b
rlabel metal1 -6 22 -6 22 5 vdd
<< end >>
