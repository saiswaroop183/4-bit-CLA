magic
tech scmos
timestamp 1638713579
<< nwell >>
rect -125 123 550 150
rect -181 4 543 31
<< ntransistor >>
rect -114 80 -112 84
rect -101 80 -99 84
rect -83 80 -81 84
rect -73 80 -71 84
rect -54 80 -52 84
rect -34 80 -32 84
rect 35 80 37 84
rect 48 80 50 84
rect 66 80 68 84
rect 76 80 78 84
rect 95 80 97 84
rect 115 80 117 84
rect 184 80 186 84
rect 197 80 199 84
rect 215 80 217 84
rect 225 80 227 84
rect 244 80 246 84
rect 264 80 266 84
rect 333 80 335 84
rect 346 80 348 84
rect 364 80 366 84
rect 374 80 376 84
rect 390 80 392 84
rect 405 80 407 84
rect 465 80 467 84
rect 478 80 480 84
rect 496 80 498 84
rect 506 80 508 84
rect 523 80 525 84
rect 537 80 539 84
rect -10 73 -8 77
rect 0 73 2 77
rect 10 73 12 77
rect 139 73 141 77
rect 149 73 151 77
rect 159 73 161 77
rect 288 73 290 77
rect 298 73 300 77
rect 308 73 310 77
rect 427 73 429 77
rect 437 73 439 77
rect 447 73 449 77
rect 38 -22 40 -18
rect 48 -22 50 -18
rect 58 -22 60 -18
rect 88 -22 90 -18
rect 98 -22 100 -18
rect 108 -22 110 -18
rect 133 -22 135 -18
rect 143 -22 145 -18
rect 153 -22 155 -18
rect 177 -22 179 -18
rect 187 -22 189 -18
rect 197 -22 199 -18
rect 215 -22 217 -18
rect 240 -22 242 -18
rect 250 -22 252 -18
rect 260 -22 262 -18
rect 278 -22 280 -18
rect 305 -22 307 -18
rect 315 -22 317 -18
rect 325 -22 327 -18
rect 336 -22 338 -18
rect 354 -22 356 -18
rect 380 -22 382 -18
rect 390 -22 392 -18
rect 400 -22 402 -18
rect 418 -22 420 -18
rect 434 -22 436 -18
rect 444 -22 446 -18
rect 454 -22 456 -18
rect 479 -22 481 -18
rect 489 -22 491 -18
rect 499 -22 501 -18
rect 510 -22 512 -18
rect 528 -22 530 -18
rect -170 -39 -168 -35
rect -157 -39 -155 -35
rect -139 -39 -137 -35
rect -129 -39 -127 -35
rect -110 -39 -108 -35
rect -90 -39 -88 -35
rect -66 -39 -64 -35
rect -53 -39 -51 -35
rect -35 -39 -33 -35
rect -25 -39 -23 -35
rect -6 -39 -4 -35
rect 14 -39 16 -35
<< ptransistor >>
rect -114 130 -112 138
rect -101 130 -99 138
rect -83 130 -81 138
rect -73 130 -71 138
rect -54 130 -52 138
rect -34 130 -32 138
rect -10 130 -8 138
rect 0 130 2 138
rect 10 130 12 138
rect 35 130 37 138
rect 48 130 50 138
rect 66 130 68 138
rect 76 130 78 138
rect 95 130 97 138
rect 115 130 117 138
rect 139 130 141 138
rect 149 130 151 138
rect 159 130 161 138
rect 184 130 186 138
rect 197 130 199 138
rect 215 130 217 138
rect 225 130 227 138
rect 244 130 246 138
rect 264 130 266 138
rect 288 130 290 138
rect 298 130 300 138
rect 308 130 310 138
rect 333 130 335 138
rect 346 130 348 138
rect 364 130 366 138
rect 374 130 376 138
rect 390 130 392 138
rect 405 130 407 138
rect 427 130 429 138
rect 437 130 439 138
rect 447 130 449 138
rect 465 130 467 138
rect 478 130 480 138
rect 496 130 498 138
rect 506 130 508 138
rect 523 130 525 138
rect 537 130 539 138
rect -170 11 -168 19
rect -157 11 -155 19
rect -139 11 -137 19
rect -129 11 -127 19
rect -110 11 -108 19
rect -90 11 -88 19
rect -66 11 -64 19
rect -53 11 -51 19
rect -35 11 -33 19
rect -25 11 -23 19
rect -6 11 -4 19
rect 14 11 16 19
rect 38 11 40 19
rect 48 11 50 19
rect 58 11 60 19
rect 88 11 90 19
rect 98 11 100 19
rect 108 11 110 19
rect 133 11 135 19
rect 143 11 145 19
rect 153 11 155 19
rect 177 11 179 19
rect 187 11 189 19
rect 197 11 199 19
rect 215 11 217 19
rect 240 11 242 19
rect 250 11 252 19
rect 260 11 262 19
rect 278 11 280 19
rect 305 11 307 19
rect 315 11 317 19
rect 325 11 327 19
rect 336 11 338 19
rect 354 11 356 19
rect 380 11 382 19
rect 390 11 392 19
rect 400 11 402 19
rect 418 11 420 19
rect 434 11 436 19
rect 444 11 446 19
rect 454 11 456 19
rect 479 11 481 19
rect 489 11 491 19
rect 499 11 501 19
rect 510 11 512 19
rect 528 11 530 19
<< ndiffusion >>
rect -115 80 -114 84
rect -112 80 -109 84
rect -105 80 -101 84
rect -99 80 -98 84
rect -84 80 -83 84
rect -81 80 -79 84
rect -75 80 -73 84
rect -71 80 -69 84
rect -65 80 -54 84
rect -52 80 -50 84
rect -46 80 -34 84
rect -32 80 -31 84
rect 34 80 35 84
rect 37 80 40 84
rect 44 80 48 84
rect 50 80 51 84
rect 65 80 66 84
rect 68 80 70 84
rect 74 80 76 84
rect 78 80 80 84
rect 84 80 95 84
rect 97 80 99 84
rect 103 80 115 84
rect 117 80 118 84
rect 183 80 184 84
rect 186 80 189 84
rect 193 80 197 84
rect 199 80 200 84
rect 214 80 215 84
rect 217 80 219 84
rect 223 80 225 84
rect 227 80 229 84
rect 233 80 244 84
rect 246 80 248 84
rect 252 80 264 84
rect 266 80 267 84
rect 332 80 333 84
rect 335 80 338 84
rect 342 80 346 84
rect 348 80 349 84
rect 363 80 364 84
rect 366 80 368 84
rect 372 80 374 84
rect 376 80 378 84
rect 382 80 390 84
rect 392 80 394 84
rect 398 80 405 84
rect 407 80 408 84
rect 464 80 465 84
rect 467 80 470 84
rect 474 80 478 84
rect 480 80 481 84
rect 495 80 496 84
rect 498 80 500 84
rect 504 80 506 84
rect 508 80 510 84
rect 514 80 523 84
rect 525 80 527 84
rect 531 80 537 84
rect 539 80 540 84
rect -11 73 -10 77
rect -8 73 0 77
rect 2 73 4 77
rect 8 73 10 77
rect 12 73 13 77
rect 138 73 139 77
rect 141 73 149 77
rect 151 73 153 77
rect 157 73 159 77
rect 161 73 162 77
rect 287 73 288 77
rect 290 73 298 77
rect 300 73 302 77
rect 306 73 308 77
rect 310 73 311 77
rect 426 73 427 77
rect 429 73 437 77
rect 439 73 441 77
rect 445 73 447 77
rect 449 73 450 77
rect 37 -22 38 -18
rect 40 -22 48 -18
rect 50 -22 52 -18
rect 56 -22 58 -18
rect 60 -22 61 -18
rect 87 -22 88 -18
rect 90 -22 92 -18
rect 96 -22 98 -18
rect 100 -22 102 -18
rect 106 -22 108 -18
rect 110 -22 111 -18
rect 132 -22 133 -18
rect 135 -22 143 -18
rect 145 -22 147 -18
rect 151 -22 153 -18
rect 155 -22 156 -18
rect 176 -22 177 -18
rect 179 -22 187 -18
rect 189 -22 197 -18
rect 199 -22 200 -18
rect 209 -22 210 -18
rect 214 -22 215 -18
rect 217 -22 218 -18
rect 239 -22 240 -18
rect 242 -22 244 -18
rect 248 -22 250 -18
rect 252 -22 254 -18
rect 258 -22 260 -18
rect 262 -22 263 -18
rect 272 -22 273 -18
rect 277 -22 278 -18
rect 280 -22 281 -18
rect 304 -22 305 -18
rect 307 -22 315 -18
rect 317 -22 325 -18
rect 327 -22 336 -18
rect 338 -22 339 -18
rect 348 -22 349 -18
rect 353 -22 354 -18
rect 356 -22 357 -18
rect 379 -22 380 -18
rect 382 -22 390 -18
rect 392 -22 400 -18
rect 402 -22 403 -18
rect 412 -22 413 -18
rect 417 -22 418 -18
rect 420 -22 421 -18
rect 433 -22 434 -18
rect 436 -22 444 -18
rect 446 -22 448 -18
rect 452 -22 454 -18
rect 456 -22 457 -18
rect 478 -22 479 -18
rect 481 -22 483 -18
rect 487 -22 489 -18
rect 491 -22 493 -18
rect 497 -22 499 -18
rect 501 -22 504 -18
rect 508 -22 510 -18
rect 512 -22 513 -18
rect 522 -22 523 -18
rect 527 -22 528 -18
rect 530 -22 531 -18
rect -171 -39 -170 -35
rect -168 -39 -165 -35
rect -161 -39 -157 -35
rect -155 -39 -154 -35
rect -140 -39 -139 -35
rect -137 -39 -135 -35
rect -131 -39 -129 -35
rect -127 -39 -125 -35
rect -121 -39 -110 -35
rect -108 -39 -106 -35
rect -102 -39 -90 -35
rect -88 -39 -87 -35
rect -67 -39 -66 -35
rect -64 -39 -61 -35
rect -57 -39 -53 -35
rect -51 -39 -50 -35
rect -36 -39 -35 -35
rect -33 -39 -31 -35
rect -27 -39 -25 -35
rect -23 -39 -21 -35
rect -17 -39 -6 -35
rect -4 -39 -2 -35
rect 2 -39 14 -35
rect 16 -39 17 -35
<< pdiffusion >>
rect -115 130 -114 138
rect -112 130 -106 138
rect -102 130 -101 138
rect -99 130 -98 138
rect -84 130 -83 138
rect -81 130 -73 138
rect -71 130 -69 138
rect -65 130 -54 138
rect -52 130 -34 138
rect -32 130 -31 138
rect -11 130 -10 138
rect -8 130 -6 138
rect -2 130 0 138
rect 2 130 4 138
rect 8 130 10 138
rect 12 130 13 138
rect 34 130 35 138
rect 37 130 43 138
rect 47 130 48 138
rect 50 130 51 138
rect 65 130 66 138
rect 68 130 76 138
rect 78 130 80 138
rect 84 130 95 138
rect 97 130 115 138
rect 117 130 118 138
rect 138 130 139 138
rect 141 130 143 138
rect 147 130 149 138
rect 151 130 153 138
rect 157 130 159 138
rect 161 130 162 138
rect 183 130 184 138
rect 186 130 192 138
rect 196 130 197 138
rect 199 130 200 138
rect 214 130 215 138
rect 217 130 225 138
rect 227 130 229 138
rect 233 130 244 138
rect 246 130 264 138
rect 266 130 267 138
rect 287 130 288 138
rect 290 130 292 138
rect 296 130 298 138
rect 300 130 302 138
rect 306 130 308 138
rect 310 130 311 138
rect 332 130 333 138
rect 335 130 341 138
rect 345 130 346 138
rect 348 130 349 138
rect 363 130 364 138
rect 366 130 374 138
rect 376 130 378 138
rect 382 130 390 138
rect 392 130 405 138
rect 407 130 408 138
rect 426 130 427 138
rect 429 130 431 138
rect 435 130 437 138
rect 439 130 441 138
rect 445 130 447 138
rect 449 130 450 138
rect 464 130 465 138
rect 467 130 473 138
rect 477 130 478 138
rect 480 130 481 138
rect 495 130 496 138
rect 498 130 506 138
rect 508 130 510 138
rect 514 130 523 138
rect 525 130 537 138
rect 539 130 540 138
rect -171 11 -170 19
rect -168 11 -162 19
rect -158 11 -157 19
rect -155 11 -154 19
rect -140 11 -139 19
rect -137 11 -129 19
rect -127 11 -125 19
rect -121 11 -110 19
rect -108 11 -90 19
rect -88 11 -87 19
rect -67 11 -66 19
rect -64 11 -58 19
rect -54 11 -53 19
rect -51 11 -50 19
rect -36 11 -35 19
rect -33 11 -25 19
rect -23 11 -21 19
rect -17 11 -6 19
rect -4 11 14 19
rect 16 11 17 19
rect 37 11 38 19
rect 40 11 42 19
rect 46 11 48 19
rect 50 11 52 19
rect 56 11 58 19
rect 60 11 61 19
rect 87 11 88 19
rect 90 11 98 19
rect 100 11 102 19
rect 106 11 108 19
rect 110 11 111 19
rect 132 11 133 19
rect 135 11 137 19
rect 141 11 143 19
rect 145 11 147 19
rect 151 11 153 19
rect 155 11 156 19
rect 176 11 177 19
rect 179 11 181 19
rect 185 11 187 19
rect 189 11 191 19
rect 195 11 197 19
rect 199 11 200 19
rect 208 11 210 19
rect 214 11 215 19
rect 217 11 218 19
rect 239 11 240 19
rect 242 11 250 19
rect 252 11 260 19
rect 262 11 263 19
rect 272 11 273 19
rect 277 11 278 19
rect 280 11 281 19
rect 304 11 305 19
rect 307 11 309 19
rect 313 11 315 19
rect 317 11 319 19
rect 323 11 325 19
rect 327 11 329 19
rect 333 11 336 19
rect 338 11 339 19
rect 348 11 349 19
rect 353 11 354 19
rect 356 11 357 19
rect 379 11 380 19
rect 382 11 384 19
rect 388 11 390 19
rect 392 11 394 19
rect 398 11 400 19
rect 402 11 403 19
rect 411 11 413 19
rect 417 11 418 19
rect 420 11 421 19
rect 433 11 434 19
rect 436 11 438 19
rect 442 11 444 19
rect 446 11 448 19
rect 452 11 454 19
rect 456 11 457 19
rect 478 11 479 19
rect 481 11 489 19
rect 491 11 499 19
rect 501 11 510 19
rect 512 11 513 19
rect 522 11 523 19
rect 527 11 528 19
rect 530 11 531 19
<< ndcontact >>
rect -119 80 -115 84
rect -109 80 -105 84
rect -98 80 -94 84
rect -88 80 -84 84
rect -79 80 -75 84
rect -69 80 -65 84
rect -50 80 -46 84
rect -31 80 -27 84
rect 30 80 34 84
rect 40 80 44 84
rect 51 80 55 84
rect 61 80 65 84
rect 70 80 74 84
rect 80 80 84 84
rect 99 80 103 84
rect 118 80 122 84
rect 179 80 183 84
rect 189 80 193 84
rect 200 80 204 84
rect 210 80 214 84
rect 219 80 223 84
rect 229 80 233 84
rect 248 80 252 84
rect 267 80 271 84
rect 328 80 332 84
rect 338 80 342 84
rect 349 80 353 84
rect 359 80 363 84
rect 368 80 372 84
rect 378 80 382 84
rect 394 80 398 84
rect 408 80 412 84
rect 460 80 464 84
rect 470 80 474 84
rect 481 80 485 84
rect 491 80 495 84
rect 500 80 504 84
rect 510 80 514 84
rect 527 80 531 84
rect 540 80 544 84
rect -15 73 -11 77
rect 4 73 8 77
rect 13 73 17 77
rect 134 73 138 77
rect 153 73 157 77
rect 162 73 166 77
rect 283 73 287 77
rect 302 73 306 77
rect 311 73 315 77
rect 422 73 426 77
rect 441 73 445 77
rect 450 73 454 77
rect 33 -22 37 -18
rect 52 -22 56 -18
rect 61 -22 65 -18
rect 83 -22 87 -18
rect 92 -22 96 -18
rect 102 -22 106 -18
rect 111 -22 115 -18
rect 128 -22 132 -18
rect 147 -22 151 -18
rect 156 -22 160 -18
rect 172 -22 176 -18
rect 200 -22 204 -18
rect 210 -22 214 -18
rect 218 -22 222 -18
rect 235 -22 239 -18
rect 244 -22 248 -18
rect 254 -22 258 -18
rect 263 -22 267 -18
rect 273 -22 277 -18
rect 281 -22 285 -18
rect 300 -22 304 -18
rect 339 -22 343 -18
rect 349 -22 353 -18
rect 357 -22 361 -18
rect 375 -22 379 -18
rect 403 -22 407 -18
rect 413 -22 417 -18
rect 421 -22 425 -18
rect 429 -22 433 -18
rect 448 -22 452 -18
rect 457 -22 461 -18
rect 474 -22 478 -18
rect 483 -22 487 -18
rect 493 -22 497 -18
rect 504 -22 508 -18
rect 513 -22 517 -18
rect 523 -22 527 -18
rect 531 -22 535 -18
rect -175 -39 -171 -35
rect -165 -39 -161 -35
rect -154 -39 -150 -35
rect -144 -39 -140 -35
rect -135 -39 -131 -35
rect -125 -39 -121 -35
rect -106 -39 -102 -35
rect -87 -39 -83 -35
rect -71 -39 -67 -35
rect -61 -39 -57 -35
rect -50 -39 -46 -35
rect -40 -39 -36 -35
rect -31 -39 -27 -35
rect -21 -39 -17 -35
rect -2 -39 2 -35
rect 17 -39 21 -35
<< pdcontact >>
rect -119 130 -115 138
rect -106 130 -102 138
rect -98 130 -94 138
rect -88 130 -84 138
rect -69 130 -65 138
rect -31 130 -27 138
rect -15 130 -11 138
rect -6 130 -2 138
rect 4 130 8 138
rect 13 130 17 138
rect 30 130 34 138
rect 43 130 47 138
rect 51 130 55 138
rect 61 130 65 138
rect 80 130 84 138
rect 118 130 122 138
rect 134 130 138 138
rect 143 130 147 138
rect 153 130 157 138
rect 162 130 166 138
rect 179 130 183 138
rect 192 130 196 138
rect 200 130 204 138
rect 210 130 214 138
rect 229 130 233 138
rect 267 130 271 138
rect 283 130 287 138
rect 292 130 296 138
rect 302 130 306 138
rect 311 130 315 138
rect 328 130 332 138
rect 341 130 345 138
rect 349 130 353 138
rect 359 130 363 138
rect 378 130 382 138
rect 408 130 412 138
rect 422 130 426 138
rect 431 130 435 138
rect 441 130 445 138
rect 450 130 454 138
rect 460 130 464 138
rect 473 130 477 138
rect 481 130 485 138
rect 491 130 495 138
rect 510 130 514 138
rect 540 130 544 138
rect -175 11 -171 19
rect -162 11 -158 19
rect -154 11 -150 19
rect -144 11 -140 19
rect -125 11 -121 19
rect -87 11 -83 19
rect -71 11 -67 19
rect -58 11 -54 19
rect -50 11 -46 19
rect -40 11 -36 19
rect -21 11 -17 19
rect 17 11 21 19
rect 33 11 37 19
rect 42 11 46 19
rect 52 11 56 19
rect 61 11 65 19
rect 83 11 87 19
rect 102 11 106 19
rect 111 11 115 19
rect 128 11 132 19
rect 137 11 141 19
rect 147 11 151 19
rect 156 11 160 19
rect 172 11 176 19
rect 181 11 185 19
rect 191 11 195 19
rect 200 11 204 19
rect 210 11 214 19
rect 218 11 222 19
rect 235 11 239 19
rect 263 11 267 19
rect 273 11 277 19
rect 281 11 285 19
rect 300 11 304 19
rect 309 11 313 19
rect 319 11 323 19
rect 329 11 333 19
rect 339 11 343 19
rect 349 11 353 19
rect 357 11 361 19
rect 375 11 379 19
rect 384 11 388 19
rect 394 11 398 19
rect 403 11 407 19
rect 413 11 417 19
rect 421 11 425 19
rect 429 11 433 19
rect 438 11 442 19
rect 448 11 452 19
rect 457 11 461 19
rect 474 11 478 19
rect 513 11 517 19
rect 523 11 527 19
rect 531 11 535 19
<< psubstratepcontact >>
rect -125 65 -121 69
rect -107 65 -103 69
rect -89 65 -85 69
rect -56 65 -52 69
rect -26 65 -22 69
rect -16 65 -12 69
rect 13 65 17 69
rect 24 65 28 69
rect 42 65 46 69
rect 60 65 64 69
rect 93 65 97 69
rect 123 65 127 69
rect 133 65 137 69
rect 162 65 166 69
rect 173 65 177 69
rect 191 65 195 69
rect 209 65 213 69
rect 242 65 246 69
rect 272 65 276 69
rect 282 65 286 69
rect 311 65 315 69
rect 322 65 326 69
rect 340 65 344 69
rect 358 65 362 69
rect 388 65 392 69
rect 413 65 417 69
rect 421 65 425 69
rect 450 65 454 69
rect 458 65 462 69
rect 472 65 476 69
rect 490 65 494 69
rect 523 65 527 69
rect 32 -30 36 -26
rect 61 -30 65 -26
rect 82 -30 86 -26
rect 111 -30 115 -26
rect 127 -30 131 -26
rect 156 -30 160 -26
rect 171 -30 175 -26
rect 200 -30 204 -26
rect 222 -30 226 -26
rect 235 -30 239 -26
rect 263 -30 267 -26
rect 285 -30 289 -26
rect 300 -30 304 -26
rect 330 -30 334 -26
rect 361 -30 365 -26
rect 374 -30 378 -26
rect 403 -30 407 -26
rect 425 -30 429 -26
rect 433 -30 437 -26
rect 457 -30 461 -26
rect 474 -30 478 -26
rect 504 -30 508 -26
rect 535 -30 539 -26
rect -163 -54 -159 -50
rect -145 -54 -141 -50
rect -112 -54 -108 -50
rect -82 -54 -78 -50
rect -61 -54 -57 -50
rect -41 -54 -37 -50
rect -8 -54 -4 -50
rect 22 -54 26 -50
<< nsubstratencontact >>
rect -121 143 -117 147
rect -96 143 -92 147
rect -88 143 -84 147
rect -69 143 -65 147
rect -28 143 -24 147
rect -15 143 -11 147
rect 14 143 18 147
rect 28 143 32 147
rect 53 143 57 147
rect 61 143 65 147
rect 80 143 84 147
rect 121 143 125 147
rect 134 143 138 147
rect 163 143 167 147
rect 177 143 181 147
rect 202 143 206 147
rect 210 143 214 147
rect 229 143 233 147
rect 270 143 274 147
rect 283 143 287 147
rect 312 143 316 147
rect 326 143 330 147
rect 351 143 355 147
rect 359 143 363 147
rect 378 143 382 147
rect 411 143 415 147
rect 422 143 426 147
rect 451 143 455 147
rect 467 143 471 147
rect 483 143 487 147
rect 491 143 495 147
rect 510 143 514 147
rect 543 143 547 147
rect -177 24 -173 28
rect -152 24 -148 28
rect -144 24 -140 28
rect -125 24 -121 28
rect -84 24 -80 28
rect -73 24 -69 28
rect -48 24 -44 28
rect -40 24 -36 28
rect -21 24 -17 28
rect 20 24 24 28
rect 33 24 37 28
rect 62 24 66 28
rect 83 24 87 28
rect 112 24 116 28
rect 128 24 132 28
rect 157 24 161 28
rect 172 24 176 28
rect 201 24 205 28
rect 220 24 224 28
rect 235 24 239 28
rect 264 24 268 28
rect 283 24 287 28
rect 300 24 304 28
rect 331 24 335 28
rect 359 24 363 28
rect 375 24 379 28
rect 404 24 408 28
rect 429 24 433 28
rect 458 24 462 28
rect 474 24 478 28
rect 505 24 509 28
rect 533 24 537 28
<< polysilicon >>
rect -114 138 -112 142
rect -101 138 -99 142
rect -83 138 -81 141
rect -73 138 -71 141
rect -54 138 -52 141
rect -34 138 -32 141
rect -10 138 -8 141
rect 0 138 2 141
rect 10 138 12 141
rect 35 138 37 142
rect 48 138 50 142
rect 66 138 68 141
rect 76 138 78 141
rect 95 138 97 141
rect 115 138 117 141
rect 139 138 141 141
rect 149 138 151 141
rect 159 138 161 141
rect 184 138 186 142
rect 197 138 199 142
rect 215 138 217 141
rect 225 138 227 141
rect 244 138 246 141
rect 264 138 266 141
rect 288 138 290 141
rect 298 138 300 141
rect 308 138 310 141
rect 333 138 335 142
rect 346 138 348 142
rect 364 138 366 141
rect 374 138 376 141
rect 390 138 392 141
rect 405 138 407 141
rect 427 138 429 141
rect 437 138 439 141
rect 447 138 449 141
rect 465 138 467 142
rect 478 138 480 142
rect 496 138 498 141
rect 506 138 508 141
rect 523 138 525 141
rect 537 138 539 141
rect -114 84 -112 130
rect -101 84 -99 130
rect -83 84 -81 130
rect -73 84 -71 130
rect -54 84 -52 130
rect -34 84 -32 130
rect -114 77 -112 80
rect -101 77 -99 80
rect -83 77 -81 80
rect -73 77 -71 80
rect -54 77 -52 80
rect -34 77 -32 80
rect -10 77 -8 130
rect 0 77 2 130
rect 10 77 12 130
rect 35 84 37 130
rect 48 84 50 130
rect 66 84 68 130
rect 76 84 78 130
rect 95 84 97 130
rect 115 84 117 130
rect 35 77 37 80
rect 48 77 50 80
rect 66 77 68 80
rect 76 77 78 80
rect 95 77 97 80
rect 115 77 117 80
rect 139 77 141 130
rect 149 77 151 130
rect 159 77 161 130
rect 184 84 186 130
rect 197 84 199 130
rect 215 84 217 130
rect 225 84 227 130
rect 244 84 246 130
rect 264 84 266 130
rect 184 77 186 80
rect 197 77 199 80
rect 215 77 217 80
rect 225 77 227 80
rect 244 77 246 80
rect 264 77 266 80
rect 288 77 290 130
rect 298 77 300 130
rect 308 77 310 130
rect 333 84 335 130
rect 346 84 348 130
rect 364 84 366 130
rect 374 84 376 130
rect 390 84 392 130
rect 405 84 407 130
rect 333 77 335 80
rect 346 77 348 80
rect 364 77 366 80
rect 374 77 376 80
rect 390 77 392 80
rect 405 77 407 80
rect 427 77 429 130
rect 437 77 439 130
rect 447 77 449 130
rect 465 84 467 130
rect 478 84 480 130
rect 496 84 498 130
rect 506 84 508 130
rect 523 84 525 130
rect 537 84 539 130
rect 465 77 467 80
rect 478 77 480 80
rect 496 77 498 80
rect 506 77 508 80
rect 523 77 525 80
rect 537 77 539 80
rect -10 70 -8 73
rect 0 70 2 73
rect 10 70 12 73
rect 139 70 141 73
rect 149 70 151 73
rect 159 70 161 73
rect 288 70 290 73
rect 298 70 300 73
rect 308 70 310 73
rect 427 70 429 73
rect 437 70 439 73
rect 447 70 449 73
rect -170 19 -168 23
rect -157 19 -155 23
rect -139 19 -137 22
rect -129 19 -127 22
rect -110 19 -108 22
rect -90 19 -88 22
rect -66 19 -64 23
rect -53 19 -51 23
rect -35 19 -33 22
rect -25 19 -23 22
rect -6 19 -4 22
rect 14 19 16 22
rect 38 19 40 35
rect 48 19 50 35
rect 58 19 60 22
rect 88 19 90 22
rect 98 19 100 35
rect 108 19 110 22
rect 133 19 135 35
rect 143 19 145 35
rect 153 19 155 22
rect 177 19 179 35
rect 187 19 189 22
rect 197 19 199 35
rect 215 19 217 22
rect 240 19 242 22
rect 250 19 252 35
rect 260 19 262 22
rect 278 19 280 22
rect 305 19 307 22
rect 315 19 317 22
rect 325 19 327 35
rect 336 19 338 35
rect 354 19 356 22
rect 380 19 382 35
rect 390 19 392 22
rect 400 19 402 35
rect 418 19 420 22
rect 434 19 436 33
rect 444 19 446 33
rect 454 19 456 22
rect 479 19 481 22
rect 489 19 491 22
rect 499 19 501 22
rect 510 19 512 36
rect 528 19 530 22
rect -170 -35 -168 11
rect -157 -35 -155 11
rect -139 -35 -137 11
rect -129 -35 -127 11
rect -110 -35 -108 11
rect -90 -35 -88 11
rect -66 -35 -64 11
rect -53 -35 -51 11
rect -35 -35 -33 11
rect -25 -35 -23 11
rect -6 -35 -4 11
rect 14 -35 16 11
rect 38 -18 40 11
rect 48 -18 50 11
rect 58 -18 60 11
rect 88 -18 90 11
rect 98 -18 100 11
rect 108 -18 110 11
rect 133 -18 135 11
rect 143 -18 145 11
rect 153 -18 155 11
rect 177 -18 179 11
rect 187 -18 189 11
rect 197 -18 199 11
rect 215 -18 217 11
rect 240 -18 242 11
rect 250 -18 252 11
rect 260 -18 262 11
rect 278 -18 280 11
rect 305 -18 307 11
rect 315 -18 317 11
rect 325 -18 327 11
rect 336 -18 338 11
rect 354 -18 356 11
rect 380 -18 382 11
rect 390 -18 392 11
rect 400 -18 402 11
rect 418 -18 420 11
rect 434 -18 436 11
rect 444 -18 446 11
rect 454 -18 456 11
rect 479 -18 481 11
rect 489 -18 491 11
rect 499 -18 501 11
rect 510 -18 512 11
rect 528 -18 530 11
rect 38 -25 40 -22
rect 48 -38 50 -22
rect 58 -25 60 -22
rect 88 -25 90 -22
rect 98 -25 100 -22
rect 108 -25 110 -22
rect 133 -25 135 -22
rect 143 -25 145 -22
rect 153 -25 155 -22
rect 177 -25 179 -22
rect 187 -39 189 -22
rect 197 -39 199 -22
rect 215 -25 217 -22
rect 240 -25 242 -22
rect 250 -25 252 -22
rect 260 -25 262 -22
rect 278 -25 280 -22
rect 305 -37 307 -22
rect 315 -37 317 -22
rect 325 -25 327 -22
rect 336 -25 338 -22
rect 354 -25 356 -22
rect 380 -25 382 -22
rect 390 -37 392 -22
rect 400 -25 402 -22
rect 418 -25 420 -22
rect 434 -25 436 -22
rect 444 -25 446 -22
rect 454 -25 456 -22
rect 479 -25 481 -22
rect 489 -25 491 -22
rect 499 -33 501 -22
rect 510 -25 512 -22
rect 528 -25 530 -22
rect -170 -42 -168 -39
rect -157 -42 -155 -39
rect -139 -42 -137 -39
rect -129 -42 -127 -39
rect -110 -42 -108 -39
rect -90 -46 -88 -39
rect -66 -42 -64 -39
rect -53 -42 -51 -39
rect -35 -42 -33 -39
rect -25 -42 -23 -39
rect -6 -42 -4 -39
rect 14 -42 16 -39
<< polycontact >>
rect -112 114 -108 118
rect -105 88 -101 92
rect -87 89 -83 93
rect -71 107 -67 111
rect -52 105 -48 109
rect -14 117 -10 121
rect -32 101 -28 105
rect -4 111 0 115
rect 6 118 10 122
rect 37 114 41 118
rect 44 88 48 92
rect 62 89 66 93
rect 78 107 82 111
rect 97 105 101 109
rect 135 117 139 121
rect 117 101 121 105
rect 145 111 149 115
rect 155 118 159 122
rect 186 114 190 118
rect 193 88 197 92
rect 211 89 215 93
rect 227 107 231 111
rect 246 105 250 109
rect 284 117 288 121
rect 266 101 270 105
rect 294 111 298 115
rect 304 118 308 122
rect 335 114 339 118
rect 342 88 346 92
rect 360 89 364 93
rect 376 107 380 111
rect 392 105 396 109
rect 423 117 427 121
rect 407 101 411 105
rect 433 111 437 115
rect 443 118 447 122
rect 467 114 471 118
rect 474 88 478 92
rect 492 89 496 93
rect 508 107 512 111
rect 525 109 529 113
rect 539 109 543 113
rect 34 31 38 35
rect 50 31 54 35
rect 100 31 104 35
rect 129 31 133 35
rect 145 31 149 35
rect 173 31 177 35
rect 199 31 203 35
rect 252 31 256 35
rect 327 31 331 35
rect 338 31 342 35
rect 376 31 380 35
rect 396 31 400 35
rect 433 33 437 37
rect 443 33 447 37
rect 506 31 510 35
rect -168 -5 -164 -1
rect -161 -31 -157 -27
rect -143 -30 -139 -26
rect -127 -12 -123 -8
rect -108 -10 -104 -6
rect -88 -10 -84 -6
rect -64 -4 -60 0
rect -57 -31 -53 -27
rect -39 -30 -35 -26
rect -23 -12 -19 -8
rect -4 -10 0 -6
rect 16 -10 20 -6
rect 54 -1 58 3
rect 84 -15 88 -11
rect 104 -9 108 -5
rect 149 -1 153 3
rect 211 -12 215 -8
rect 236 -2 240 2
rect 256 -2 260 2
rect 274 -12 278 -8
rect 350 -12 354 -8
rect 414 -12 418 -8
rect 450 -1 454 3
rect 475 -15 479 -11
rect 485 -2 489 2
rect 524 -12 528 -8
rect 50 -37 54 -33
rect 183 -37 187 -33
rect 199 -37 203 -33
rect 301 -37 305 -33
rect 311 -37 315 -33
rect 386 -37 390 -33
rect 498 -37 502 -33
rect -88 -46 -84 -42
<< metal1 >>
rect -144 143 -121 147
rect -117 143 -96 147
rect -92 143 -88 147
rect -84 143 -69 147
rect -65 143 -28 147
rect -24 143 -15 147
rect -11 143 14 147
rect 18 143 28 147
rect 32 143 53 147
rect 57 143 61 147
rect 65 143 80 147
rect 84 143 121 147
rect 125 143 134 147
rect 138 143 163 147
rect 167 143 177 147
rect 181 143 202 147
rect 206 143 210 147
rect 214 143 229 147
rect 233 143 270 147
rect 274 143 283 147
rect 287 143 312 147
rect 316 143 326 147
rect 330 143 351 147
rect 355 143 359 147
rect 363 143 378 147
rect 382 143 411 147
rect 415 143 422 147
rect 426 143 451 147
rect 455 143 467 147
rect 471 143 483 147
rect 487 143 491 147
rect 495 143 510 147
rect 514 143 543 147
rect -144 28 -140 143
rect -106 138 -102 143
rect -69 138 -65 143
rect -15 138 -11 143
rect 4 138 8 143
rect 43 138 47 143
rect 80 138 84 143
rect 134 138 138 143
rect 153 138 157 143
rect 192 138 196 143
rect 229 138 233 143
rect 283 138 287 143
rect 302 138 306 143
rect 341 138 345 143
rect 378 138 382 143
rect 422 138 426 143
rect 441 138 445 143
rect 473 138 477 143
rect 510 138 514 143
rect -119 90 -115 130
rect -108 114 -107 118
rect -98 93 -94 130
rect -88 121 -84 130
rect -31 121 -27 130
rect -6 122 -2 130
rect -88 116 -27 121
rect -79 112 -75 116
rect -18 117 -14 120
rect -6 118 6 122
rect -67 107 -66 111
rect -122 86 -115 90
rect -106 88 -105 92
rect -98 89 -87 93
rect -119 84 -115 86
rect -98 84 -94 89
rect -79 84 -75 107
rect -48 105 -44 109
rect -7 105 -4 115
rect -28 101 -24 105
rect -19 101 -4 105
rect -69 87 -27 91
rect -69 84 -65 87
rect -31 84 -27 87
rect 4 84 8 118
rect -109 69 -105 80
rect -88 76 -84 80
rect -69 76 -65 80
rect -88 72 -65 76
rect -15 80 8 84
rect 13 84 17 130
rect 30 90 34 130
rect 41 114 42 118
rect 51 93 55 130
rect 61 121 65 130
rect 118 121 122 130
rect 143 122 147 130
rect 61 116 122 121
rect 70 112 74 116
rect 131 117 135 120
rect 143 118 155 122
rect 82 107 83 111
rect 27 86 34 90
rect 43 88 44 92
rect 51 89 62 93
rect 30 84 34 86
rect 51 84 55 89
rect 70 84 74 107
rect 101 105 105 109
rect 142 105 145 115
rect 121 101 125 105
rect 130 101 145 105
rect -50 69 -46 80
rect -15 77 -11 80
rect 80 87 122 91
rect 80 84 84 87
rect 118 84 122 87
rect 153 84 157 118
rect 13 77 17 79
rect 4 69 8 73
rect 40 69 44 80
rect 61 76 65 80
rect 80 76 84 80
rect 61 72 84 76
rect 134 80 157 84
rect 162 86 166 130
rect 179 95 183 130
rect 190 114 191 118
rect 176 91 183 95
rect 200 93 204 130
rect 210 121 214 130
rect 267 121 271 130
rect 292 122 296 130
rect 210 116 271 121
rect 219 112 223 116
rect 280 117 284 120
rect 292 118 304 122
rect 231 107 232 111
rect 179 84 183 91
rect 192 88 193 92
rect 200 89 211 93
rect 200 84 204 89
rect 219 84 223 107
rect 250 105 254 109
rect 291 105 294 115
rect 270 101 274 105
rect 279 101 294 105
rect 99 69 103 80
rect 134 77 138 80
rect 162 77 166 81
rect 229 87 271 91
rect 229 84 233 87
rect 267 84 271 87
rect 302 84 306 118
rect 153 69 157 73
rect 189 69 193 80
rect 210 76 214 80
rect 229 76 233 80
rect 210 72 233 76
rect 283 80 306 84
rect 311 113 315 130
rect 311 110 317 113
rect 311 85 315 110
rect 328 95 332 130
rect 339 114 340 118
rect 325 91 332 95
rect 349 93 353 130
rect 359 121 363 130
rect 408 121 412 130
rect 431 122 435 130
rect 359 116 412 121
rect 368 112 372 116
rect 421 117 423 120
rect 431 118 443 122
rect 380 107 381 111
rect 328 84 332 91
rect 341 88 342 92
rect 349 89 360 93
rect 349 84 353 89
rect 368 84 372 107
rect 396 105 399 109
rect 430 105 433 115
rect 411 101 415 105
rect 420 101 433 105
rect 378 87 412 91
rect 378 84 382 87
rect 408 84 412 87
rect 441 84 445 118
rect 248 69 252 80
rect 283 77 287 80
rect 311 77 315 80
rect 302 69 306 73
rect 338 69 342 80
rect 359 76 363 80
rect 378 76 382 80
rect 359 72 382 76
rect 422 80 445 84
rect 450 82 454 130
rect 460 104 464 130
rect 471 114 472 118
rect 460 84 464 99
rect 481 93 485 130
rect 491 121 495 130
rect 540 121 544 130
rect 491 116 544 121
rect 500 112 504 116
rect 512 107 513 111
rect 529 109 531 113
rect 543 109 544 113
rect 473 88 474 92
rect 481 89 492 93
rect 481 84 485 89
rect 500 84 504 107
rect 394 69 398 80
rect 422 77 426 80
rect 510 87 544 91
rect 510 84 514 87
rect 540 84 544 87
rect 441 69 445 73
rect 470 69 474 80
rect 491 76 495 80
rect 510 76 514 80
rect 491 72 514 76
rect 527 69 531 80
rect -121 65 -107 69
rect -103 65 -89 69
rect -85 65 -56 69
rect -52 65 -26 69
rect -22 65 -16 69
rect -12 65 13 69
rect 17 65 24 69
rect 28 65 42 69
rect 46 65 60 69
rect 64 65 93 69
rect 97 65 123 69
rect 127 65 133 69
rect 137 65 162 69
rect 166 65 173 69
rect 177 65 191 69
rect 195 65 209 69
rect 213 65 242 69
rect 246 65 272 69
rect 276 65 282 69
rect 286 65 311 69
rect 315 65 322 69
rect 326 65 340 69
rect 344 65 358 69
rect 362 65 388 69
rect 392 65 413 69
rect 417 65 421 69
rect 425 65 450 69
rect 454 65 458 69
rect 462 65 472 69
rect 476 65 490 69
rect 494 65 523 69
rect 527 65 543 69
rect 13 35 18 41
rect 57 35 60 56
rect 186 54 189 57
rect 111 35 116 49
rect 146 51 203 54
rect 146 35 149 51
rect 174 35 177 41
rect 200 35 203 51
rect 312 38 315 57
rect 358 46 361 57
rect 358 41 360 46
rect 13 31 34 35
rect 54 31 60 35
rect 104 31 129 35
rect 256 33 312 34
rect 328 35 331 41
rect 256 31 317 33
rect 358 34 361 41
rect 396 35 399 50
rect 424 43 447 46
rect 342 31 376 34
rect 444 37 447 43
rect 424 34 433 37
rect 437 34 439 37
rect 503 31 506 34
rect -173 24 -152 28
rect -148 24 -144 28
rect -140 24 -125 28
rect -121 24 -84 28
rect -80 24 -73 28
rect -69 24 -48 28
rect -44 24 -40 28
rect -36 24 -21 28
rect -17 24 20 28
rect 24 24 33 28
rect 37 24 62 28
rect 66 24 83 28
rect 87 24 112 28
rect 116 24 128 28
rect 132 24 157 28
rect 161 24 172 28
rect 176 24 201 28
rect 205 24 220 28
rect 224 24 235 28
rect 239 24 264 28
rect 268 24 283 28
rect 287 24 300 28
rect 304 24 331 28
rect 335 24 359 28
rect 363 24 375 28
rect 379 24 404 28
rect 408 24 429 28
rect 433 24 458 28
rect 462 24 474 28
rect 478 24 505 28
rect 509 24 533 28
rect -162 19 -158 24
rect -125 19 -121 24
rect -58 19 -54 24
rect -21 19 -17 24
rect 33 19 37 24
rect 52 19 56 24
rect 102 19 106 24
rect 128 19 132 24
rect 147 19 151 24
rect 172 19 176 24
rect 191 19 195 24
rect 210 19 214 24
rect 235 19 239 24
rect 273 19 277 24
rect 300 19 304 24
rect 319 19 323 24
rect 339 19 343 24
rect -175 -15 -171 11
rect -164 -5 -163 -1
rect -175 -35 -171 -20
rect -154 -26 -150 11
rect -144 2 -140 11
rect -87 2 -83 11
rect -144 -3 -83 2
rect -135 -7 -131 -3
rect -123 -12 -122 -8
rect -104 -10 -100 -6
rect -84 -10 -80 -6
rect -162 -31 -161 -27
rect -154 -30 -143 -26
rect -154 -35 -150 -30
rect -135 -35 -131 -12
rect -71 -15 -67 11
rect -60 -4 -59 0
rect -125 -32 -83 -28
rect -125 -35 -121 -32
rect -87 -35 -83 -32
rect -165 -50 -161 -39
rect -144 -43 -140 -39
rect -125 -43 -121 -39
rect -144 -47 -121 -43
rect -71 -35 -67 -20
rect -50 -26 -46 11
rect -40 2 -36 11
rect 17 2 21 11
rect -40 -3 21 2
rect 42 3 46 11
rect 42 -1 54 3
rect -31 -7 -27 -3
rect -19 -12 -18 -8
rect 0 -10 4 -7
rect 20 -10 24 -6
rect 52 -11 56 -1
rect -58 -31 -57 -27
rect -50 -30 -39 -26
rect -50 -35 -46 -30
rect -31 -35 -27 -12
rect 33 -15 56 -11
rect 61 -12 65 11
rect 349 19 353 24
rect 375 19 379 24
rect 394 19 398 24
rect 413 19 417 24
rect 429 19 433 24
rect 448 19 452 24
rect 474 19 478 24
rect 523 19 527 24
rect 83 -5 87 11
rect 83 -8 104 -5
rect 61 -15 84 -12
rect 33 -18 37 -15
rect 61 -18 65 -15
rect 92 -18 96 -8
rect 111 -6 115 11
rect 137 3 141 11
rect 137 -1 149 3
rect 147 -11 151 -1
rect 111 -18 115 -11
rect 128 -15 151 -11
rect 156 -10 160 11
rect 181 3 185 11
rect 200 3 204 11
rect 181 -1 204 3
rect 200 -8 204 -1
rect 218 -6 222 11
rect 230 -2 236 1
rect 254 -2 256 2
rect 254 -6 257 -2
rect 156 -15 159 -10
rect 200 -12 211 -8
rect 218 -9 257 -6
rect 263 -8 267 11
rect 128 -18 132 -15
rect 156 -18 160 -15
rect 200 -18 204 -12
rect 218 -18 222 -9
rect 263 -12 274 -8
rect 244 -15 267 -12
rect 244 -18 248 -15
rect 263 -18 267 -15
rect 281 -18 285 11
rect 309 -1 313 11
rect 329 -1 333 11
rect 309 -4 343 -1
rect 339 -8 343 -4
rect 339 -12 350 -8
rect 339 -18 343 -12
rect 357 -18 361 11
rect 384 3 388 11
rect 403 3 407 11
rect 384 -1 407 3
rect 403 -8 407 -1
rect 403 -12 414 -8
rect 421 -9 425 11
rect 438 3 442 11
rect 438 -1 450 3
rect 403 -18 407 -12
rect 448 -11 452 -1
rect 421 -18 425 -14
rect 429 -15 452 -11
rect 457 -11 461 11
rect 476 -2 485 1
rect 513 -8 517 11
rect 531 -2 535 11
rect 531 -6 537 -2
rect 457 -15 475 -11
rect 513 -12 524 -8
rect 483 -15 517 -12
rect 429 -18 433 -15
rect 457 -18 461 -15
rect 483 -18 487 -15
rect 504 -18 508 -15
rect 531 -18 535 -6
rect 52 -26 56 -22
rect 83 -26 87 -22
rect 102 -26 106 -22
rect 147 -26 151 -22
rect 172 -26 176 -22
rect 210 -26 214 -22
rect 235 -26 239 -22
rect 254 -26 258 -22
rect 273 -26 277 -22
rect 300 -26 304 -22
rect 349 -26 353 -22
rect 375 -26 379 -22
rect 413 -26 417 -22
rect 448 -26 452 -22
rect 474 -26 478 -22
rect 493 -26 497 -22
rect 513 -26 517 -22
rect 523 -26 527 -22
rect 540 -26 543 65
rect -21 -32 21 -28
rect -21 -35 -17 -32
rect 17 -35 21 -32
rect -106 -50 -102 -39
rect -84 -46 -82 -42
rect -61 -50 -57 -39
rect -40 -43 -36 -39
rect -21 -43 -17 -39
rect -40 -47 -17 -43
rect 36 -30 61 -26
rect 65 -30 82 -26
rect 86 -30 111 -26
rect 115 -30 127 -26
rect 131 -30 156 -26
rect 160 -30 171 -26
rect 175 -30 200 -26
rect 204 -30 222 -26
rect 226 -30 235 -26
rect 239 -30 263 -26
rect 267 -30 285 -26
rect 289 -30 300 -26
rect 304 -30 330 -26
rect 334 -30 361 -26
rect 365 -30 374 -26
rect 378 -30 403 -26
rect 407 -30 425 -26
rect 429 -30 433 -26
rect 437 -30 457 -26
rect 461 -30 474 -26
rect 478 -30 504 -26
rect 508 -30 535 -26
rect 539 -30 543 -26
rect -2 -50 2 -39
rect 32 -50 36 -30
rect 54 -37 183 -34
rect 203 -34 301 -33
rect 203 -36 293 -34
rect 59 -42 64 -37
rect 184 -42 187 -37
rect 298 -36 301 -34
rect 312 -42 315 -37
rect 383 -37 386 -34
rect 495 -37 498 -34
rect 184 -45 315 -42
rect -165 -54 -163 -50
rect -159 -54 -145 -50
rect -141 -54 -112 -50
rect -108 -54 -82 -50
rect -78 -54 -61 -50
rect -57 -54 -41 -50
rect -37 -54 -8 -50
rect -4 -54 22 -50
rect 26 -54 36 -50
<< m2contact >>
rect -127 86 -122 91
rect -107 114 -102 119
rect -23 115 -18 120
rect -79 107 -74 112
rect -66 107 -61 112
rect -111 88 -106 93
rect -44 104 -39 109
rect -24 100 -19 105
rect 22 86 27 91
rect 42 114 47 119
rect 126 115 131 120
rect 70 107 75 112
rect 83 107 88 112
rect 38 88 43 93
rect 105 104 110 109
rect 125 100 130 105
rect 13 79 18 84
rect 171 91 176 96
rect 191 114 196 119
rect 275 115 280 120
rect 219 107 224 112
rect 232 107 237 112
rect 162 81 167 86
rect 187 88 192 93
rect 254 104 259 109
rect 274 100 279 105
rect 320 91 325 96
rect 340 114 345 119
rect 416 115 421 120
rect 368 107 373 112
rect 381 107 386 112
rect 311 80 316 85
rect 336 88 341 93
rect 399 104 404 109
rect 415 100 420 105
rect 472 114 477 119
rect 460 99 465 104
rect 500 107 505 112
rect 513 107 518 112
rect 531 108 536 113
rect 544 108 549 113
rect 450 77 455 82
rect 56 56 61 61
rect 186 57 191 62
rect 311 57 316 62
rect 357 57 362 62
rect 111 49 116 54
rect 174 41 179 46
rect 396 50 401 55
rect 327 41 332 46
rect 360 41 365 46
rect 312 33 317 38
rect 419 42 424 47
rect 419 33 424 38
rect 498 31 503 36
rect -163 -5 -158 0
rect -175 -20 -170 -15
rect -135 -12 -130 -7
rect -122 -12 -117 -7
rect -100 -11 -95 -6
rect -80 -11 -75 -6
rect -167 -31 -162 -26
rect -59 -4 -54 1
rect -72 -20 -67 -15
rect -31 -12 -26 -7
rect -18 -12 -13 -7
rect 4 -11 9 -6
rect 24 -11 29 -6
rect -63 -31 -58 -26
rect 111 -11 116 -6
rect 225 -2 230 3
rect 159 -15 164 -10
rect 361 -3 366 2
rect 421 -14 426 -9
rect 471 -3 476 2
rect -82 -47 -77 -42
rect 59 -47 64 -42
rect 293 -39 298 -34
rect 378 -38 383 -33
rect 490 -39 495 -34
<< metal2 >>
rect -129 116 -107 119
rect -102 116 -23 119
rect -63 115 -23 116
rect 20 116 42 119
rect -63 112 -59 115
rect 47 116 126 119
rect 86 115 126 116
rect 169 116 191 119
rect 86 112 90 115
rect 196 116 275 119
rect 235 115 275 116
rect 318 116 340 119
rect 235 112 239 115
rect 345 116 416 119
rect 384 115 416 116
rect 460 116 472 119
rect 384 112 388 115
rect 477 116 520 119
rect 516 112 520 116
rect -129 107 -79 110
rect -61 107 -59 112
rect 62 107 70 110
rect 88 107 90 112
rect -44 103 -40 104
rect -126 100 -40 103
rect 211 107 219 110
rect 237 107 239 112
rect 105 100 109 104
rect -126 91 -123 100
rect -24 91 -21 100
rect 23 97 109 100
rect 361 108 368 111
rect 386 107 388 112
rect 254 103 258 104
rect 172 100 258 103
rect 398 104 399 107
rect 491 107 500 110
rect 518 107 520 112
rect 398 103 402 104
rect 321 100 402 103
rect 23 91 26 97
rect -106 88 -21 91
rect -102 76 -99 88
rect 125 91 128 100
rect 172 96 175 100
rect 43 88 128 91
rect 274 91 277 100
rect 321 96 324 100
rect 192 88 277 91
rect 415 91 418 100
rect 531 103 534 108
rect 465 100 534 103
rect 341 88 418 91
rect 545 91 548 108
rect 473 88 548 91
rect -129 73 -99 76
rect -163 0 -159 41
rect -58 1 -55 57
rect 13 46 18 79
rect 47 76 50 88
rect 26 73 50 76
rect 57 61 60 71
rect 163 53 166 81
rect 196 76 199 88
rect 175 73 199 76
rect 312 62 315 80
rect 345 76 348 88
rect 357 76 360 77
rect 324 73 348 76
rect 357 62 360 71
rect 191 58 195 61
rect 116 50 396 53
rect 18 42 174 45
rect 179 42 327 45
rect 365 43 419 46
rect 317 34 419 37
rect 451 34 454 77
rect 451 31 498 34
rect -158 -3 -115 0
rect -119 -7 -115 -3
rect -54 -3 -11 0
rect -143 -12 -135 -9
rect -117 -12 -115 -7
rect -15 -7 -11 -3
rect 160 -2 225 1
rect -100 -16 -97 -11
rect -170 -19 -97 -16
rect -80 -28 -77 -11
rect -40 -12 -31 -9
rect -13 -12 -11 -7
rect 29 -10 111 -7
rect 160 -10 163 -2
rect 366 -3 471 0
rect 5 -16 8 -11
rect -67 -19 8 -16
rect -162 -31 -77 -28
rect 24 -28 27 -11
rect -58 -31 27 -28
rect 298 -37 378 -34
rect 422 -34 425 -14
rect 422 -37 490 -34
rect -77 -46 59 -43
<< m3contact >>
rect 455 115 460 120
rect 57 106 62 111
rect 206 107 211 112
rect 356 107 361 112
rect -59 57 -54 62
rect -164 41 -158 46
rect 56 71 61 76
rect 356 71 361 76
rect 195 57 200 62
<< m123contact >>
rect 468 88 473 93
rect 13 41 18 46
rect 285 -7 290 -2
<< metal3 >>
rect 205 112 212 113
rect 56 111 63 112
rect 56 106 57 111
rect 62 106 63 111
rect 205 107 206 112
rect 211 107 212 112
rect 456 111 459 115
rect 361 108 459 111
rect 205 106 212 107
rect 56 105 63 106
rect 57 76 60 105
rect 194 62 201 63
rect 194 61 195 62
rect -54 58 195 61
rect 194 57 195 58
rect 200 61 201 62
rect 209 61 212 106
rect 357 76 360 107
rect 200 58 212 61
rect 200 57 201 58
rect 194 56 201 57
rect -158 42 13 45
rect 469 -3 472 88
rect 290 -6 472 -3
<< labels >>
rlabel metal2 -128 73 -128 76 3 a0
rlabel metal2 -129 116 -129 119 3 b0
rlabel metal1 99 145 99 145 5 vdd
rlabel metal1 79 67 79 67 1 gnd
rlabel metal2 20 116 20 119 1 b1
rlabel metal2 169 116 169 119 1 b2
rlabel metal1 317 110 317 113 1 g2
rlabel metal2 318 116 318 119 1 b3
rlabel metal2 27 73 27 76 1 a1
rlabel metal2 176 73 176 76 1 a2
rlabel metal2 325 73 325 76 1 a3
rlabel metal2 -128 107 -128 110 3 sum0
rlabel metal1 15 93 15 98 1 c1
rlabel m2contact 358 58 361 58 1 p3
rlabel m2contact 113 54 116 54 6 g1
rlabel metal2 -40 -12 -40 -9 1 sum2
rlabel metal2 -143 -12 -143 -9 1 sum1
rlabel metal1 282 -5 284 -5 1 c3
rlabel metal1 113 -3 115 -3 1 c2
rlabel metal1 537 -6 537 -2 1 c4
rlabel space 311 55 315 55 6 g2
rlabel metal2 491 107 491 110 1 sum3
<< end >>
