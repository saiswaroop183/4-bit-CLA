magic
tech scmos
timestamp 1637320003
<< nwell >>
rect -27 0 18 27
<< ntransistor >>
rect -16 -26 -14 -22
rect -6 -26 -4 -22
rect 4 -26 6 -22
<< ptransistor >>
rect -16 7 -14 15
rect -6 7 -4 15
rect 4 7 6 15
<< ndiffusion >>
rect -17 -26 -16 -22
rect -14 -26 -6 -22
rect -4 -26 -2 -22
rect 2 -26 4 -22
rect 6 -26 7 -22
<< pdiffusion >>
rect -17 7 -16 15
rect -14 7 -12 15
rect -8 7 -6 15
rect -4 7 -2 15
rect 2 7 4 15
rect 6 7 7 15
<< ndcontact >>
rect -21 -26 -17 -22
rect -2 -26 2 -22
rect 7 -26 11 -22
<< pdcontact >>
rect -21 7 -17 15
rect -12 7 -8 15
rect -2 7 2 15
rect 7 7 11 15
<< psubstratepcontact >>
rect -22 -34 -18 -30
rect 7 -34 11 -30
<< nsubstratencontact >>
rect -21 20 -17 24
rect 8 20 12 24
<< polysilicon >>
rect -16 15 -14 18
rect -6 15 -4 18
rect 4 15 6 18
rect -16 -22 -14 7
rect -6 -22 -4 7
rect 4 -22 6 7
rect -16 -29 -14 -26
rect -6 -29 -4 -26
rect 4 -29 6 -26
<< polycontact >>
rect -20 -12 -16 -8
rect -10 -12 -6 -8
rect 0 -5 4 -1
<< metal1 >>
rect -17 20 8 24
rect -21 15 -17 20
rect -2 15 2 20
rect -12 -1 -8 7
rect -12 -5 0 -1
rect -22 -12 -20 -8
rect -12 -12 -10 -8
rect -2 -15 2 -5
rect -21 -19 2 -15
rect 7 -9 11 7
rect 7 -13 13 -9
rect -21 -22 -17 -19
rect 7 -22 11 -13
rect -2 -30 2 -26
rect -18 -34 7 -30
<< labels >>
rlabel metal1 -6 22 -6 22 5 vdd
rlabel metal1 -5 -32 -5 -32 1 gnd
rlabel metal1 13 -13 13 -9 7 g
rlabel metal1 -22 -12 -22 -8 3 a
rlabel metal1 -12 -12 -12 -8 1 b
<< end >>
